-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 13 2025 20:50:07

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__49949\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49938\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49892\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49817\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49757\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49670\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49646\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49622\ : std_logic;
signal \N__49621\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49607\ : std_logic;
signal \N__49604\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49556\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49529\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49511\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49400\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49391\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49385\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49370\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49310\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49284\ : std_logic;
signal \N__49283\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49279\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49276\ : std_logic;
signal \N__49275\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49256\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49199\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49175\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49171\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49072\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48983\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48912\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48818\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48630\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48470\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48380\ : std_logic;
signal \N__48379\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47186\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47168\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47159\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46612\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45325\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45109\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44855\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44825\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44377\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44027\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43307\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42410\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42386\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42332\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41906\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41759\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \N_34_i_i\ : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_168_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_166\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_166_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_162\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \current_shift_inst.PI_CTRL.N_167\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_3_10_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \current_shift_inst.PI_CTRL.N_53\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \delay_measurement_inst.N_34\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_\ : std_logic;
signal \delay_measurement_inst.N_32\ : std_logic;
signal \delay_measurement_inst.N_35\ : std_logic;
signal \delay_measurement_inst.N_43\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_enablelt3_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_71\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal s4_phy_c : std_logic;
signal \delay_measurement_inst.N_31\ : std_logic;
signal \delay_measurement_inst.N_40\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt14_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0\ : std_logic;
signal \delay_measurement_inst.un1_elapsed_time_hc_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\ : std_logic;
signal \delay_measurement_inst.N_30_cascade_\ : std_logic;
signal \delay_measurement_inst.N_37\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_302_i\ : std_logic;
signal \delay_measurement_inst.N_36\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_72\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt30_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt14_0\ : std_logic;
signal \delay_measurement_inst.N_41\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_302_i_g\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.N_52\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.prev_hc_sigZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_16\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \bfn_10_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_30\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto15\ : std_logic;
signal \delay_measurement_inst.N_39_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_27\ : std_logic;
signal s3_phy_c : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_21\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_8\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_0_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto9\ : std_logic;
signal \delay_measurement_inst.N_33_cascade_\ : std_logic;
signal \delay_measurement_inst.N_38\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_303_i\ : std_logic;
signal \delay_measurement_inst.N_28\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal measured_delay_hc_25 : std_logic;
signal measured_delay_hc_24 : std_logic;
signal measured_delay_hc_26 : std_logic;
signal measured_delay_hc_23 : std_logic;
signal measured_delay_hc_28 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.N_51\ : std_logic;
signal measured_delay_hc_27 : std_logic;
signal \delay_measurement_inst.N_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_304_i\ : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal delay_tr_d2 : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.prev_tr_sigZ0\ : std_logic;
signal \delay_measurement_inst.N_59\ : std_logic;
signal \delay_measurement_inst.N_270\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal measured_delay_hc_14 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal measured_delay_hc_19 : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal measured_delay_hc_17 : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3\ : std_logic;
signal measured_delay_hc_20 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.N_29_cascade_\ : std_logic;
signal measured_delay_hc_6 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6\ : std_logic;
signal measured_delay_hc_21 : std_logic;
signal \delay_measurement_inst.N_42\ : std_logic;
signal measured_delay_hc_18 : std_logic;
signal \delay_measurement_inst.N_26\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \delay_measurement_inst.N_27\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.N_53\ : std_logic;
signal measured_delay_hc_29 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3\ : std_logic;
signal \delay_measurement_inst.N_54\ : std_logic;
signal measured_delay_hc_30 : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal delay_hc_d2 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\ : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7\ : std_logic;
signal \delay_measurement_inst.N_299\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal measured_delay_hc_4 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal measured_delay_hc_5 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal measured_delay_hc_16 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal measured_delay_hc_1 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_start\ : std_logic;
signal measured_delay_hc_3 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal measured_delay_hc_7 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal measured_delay_hc_8 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal measured_delay_hc_0 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal measured_delay_hc_13 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal measured_delay_hc_15 : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt30\ : std_logic;
signal measured_delay_hc_2 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal measured_delay_hc_12 : std_logic;
signal measured_delay_hc_11 : std_logic;
signal measured_delay_hc_9 : std_logic;
signal measured_delay_hc_10 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.un1_elapsed_time_hc\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lt31_0\ : std_logic;
signal measured_delay_hc_22 : std_logic;
signal state_3 : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_181_i\ : std_logic;
signal s2_phy_c : std_logic;
signal \phase_controller_inst2.stoper_tr.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal measured_delay_tr_5 : std_logic;
signal measured_delay_tr_3 : std_logic;
signal \phase_controller_inst1.stoper_tr.N_248\ : std_logic;
signal measured_delay_tr_1 : std_logic;
signal measured_delay_tr_11 : std_logic;
signal measured_delay_tr_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\ : std_logic;
signal measured_delay_tr_6 : std_logic;
signal measured_delay_tr_2 : std_logic;
signal \phase_controller_inst1.stoper_tr.N_55\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal red_c_i : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_RNO_0_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal measured_delay_hc_31 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_15_2_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \bfn_15_3_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \bfn_15_4_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_290\ : std_logic;
signal \delay_measurement_inst.N_325\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal measured_delay_tr_10 : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\ : std_logic;
signal measured_delay_tr_4 : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\ : std_logic;
signal measured_delay_tr_19 : std_logic;
signal measured_delay_tr_12 : std_logic;
signal measured_delay_tr_14 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\ : std_logic;
signal measured_delay_tr_13 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\ : std_logic;
signal measured_delay_tr_15 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal measured_delay_tr_17 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal measured_delay_tr_18 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal measured_delay_tr_7 : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i\ : std_logic;
signal \delay_measurement_inst.N_267\ : std_logic;
signal measured_delay_tr_8 : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.N_1318_i\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_1_axb_11\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_15_27_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_15_28_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_181_i_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\ : std_logic;
signal \delay_measurement_inst.N_265\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_287_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal \bfn_16_7_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \bfn_16_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un4_control_input_0_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal measured_delay_tr_16 : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_305_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_304_i_g\ : std_logic;
signal start_stop_c : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \current_shift_inst.timer_s1.N_180_i_g\ : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21250\&\N__21176\&\N__21248\&\N__21175\&\N__21249\&\N__21174\&\N__21251\&\N__21171\&\N__21244\&\N__21170\&\N__21245\&\N__21172\&\N__21246\&\N__21173\&\N__21247\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__46030\&\N__46027\&'0'&'0'&'0'&\N__46025\&\N__46029\&\N__46026\&\N__46028\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21261\&\N__21264\&\N__21262\&\N__21265\&\N__21263\&\N__20319\&\N__20265\&\N__21033\&\N__20295\&\N__21006\&\N__20209\&\N__20249\&\N__19976\&\N__19991\&\N__20006\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__45896\&\N__45893\&'0'&'0'&'0'&\N__45891\&\N__45895\&\N__45892\&\N__45894\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__24662\,
            RESETB => \N__35913\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__46031\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__46024\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__45857\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__45890\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__49947\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49949\,
            DIN => \N__49948\,
            DOUT => \N__49947\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49949\,
            PADOUT => \N__49948\,
            PADIN => \N__49947\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49938\,
            DIN => \N__49937\,
            DOUT => \N__49936\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49938\,
            PADOUT => \N__49937\,
            PADIN => \N__49936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49929\,
            DIN => \N__49928\,
            DOUT => \N__49927\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49929\,
            PADOUT => \N__49928\,
            PADIN => \N__49927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49920\,
            DIN => \N__49919\,
            DOUT => \N__49918\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49920\,
            PADOUT => \N__49919\,
            PADIN => \N__49918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21893\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49911\,
            DIN => \N__49910\,
            DOUT => \N__49909\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49911\,
            PADOUT => \N__49910\,
            PADIN => \N__49909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49902\,
            DIN => \N__49901\,
            DOUT => \N__49900\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49902\,
            PADOUT => \N__49901\,
            PADIN => \N__49900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34520\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49893\,
            DIN => \N__49892\,
            DOUT => \N__49891\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49893\,
            PADOUT => \N__49892\,
            PADIN => \N__49891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49884\,
            DIN => \N__49883\,
            DOUT => \N__49882\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49884\,
            PADOUT => \N__49883\,
            PADIN => \N__49882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49875\,
            DIN => \N__49874\,
            DOUT => \N__49873\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49875\,
            PADOUT => \N__49874\,
            PADIN => \N__49873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49866\,
            DIN => \N__49865\,
            DOUT => \N__49864\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49866\,
            PADOUT => \N__49865\,
            PADIN => \N__49864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34574\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49857\,
            DIN => \N__49856\,
            DOUT => \N__49855\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49857\,
            PADOUT => \N__49856\,
            PADIN => \N__49855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23249\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49848\,
            DIN => \N__49847\,
            DOUT => \N__49846\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49848\,
            PADOUT => \N__49847\,
            PADIN => \N__49846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49839\,
            DIN => \N__49838\,
            DOUT => \N__49837\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49839\,
            PADOUT => \N__49838\,
            PADIN => \N__49837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11854\ : InMux
    port map (
            O => \N__49820\,
            I => \N__49817\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__49817\,
            I => \N__49814\
        );

    \I__11852\ : Odrv12
    port map (
            O => \N__49814\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__11851\ : InMux
    port map (
            O => \N__49811\,
            I => \N__49808\
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__49808\,
            I => \N__49805\
        );

    \I__11849\ : Odrv12
    port map (
            O => \N__49805\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__11848\ : InMux
    port map (
            O => \N__49802\,
            I => \N__49799\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__49799\,
            I => \N__49796\
        );

    \I__11846\ : Span4Mux_h
    port map (
            O => \N__49796\,
            I => \N__49793\
        );

    \I__11845\ : Odrv4
    port map (
            O => \N__49793\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__11844\ : InMux
    port map (
            O => \N__49790\,
            I => \N__49787\
        );

    \I__11843\ : LocalMux
    port map (
            O => \N__49787\,
            I => \N__49772\
        );

    \I__11842\ : InMux
    port map (
            O => \N__49786\,
            I => \N__49767\
        );

    \I__11841\ : InMux
    port map (
            O => \N__49785\,
            I => \N__49767\
        );

    \I__11840\ : InMux
    port map (
            O => \N__49784\,
            I => \N__49758\
        );

    \I__11839\ : InMux
    port map (
            O => \N__49783\,
            I => \N__49729\
        );

    \I__11838\ : InMux
    port map (
            O => \N__49782\,
            I => \N__49716\
        );

    \I__11837\ : InMux
    port map (
            O => \N__49781\,
            I => \N__49716\
        );

    \I__11836\ : InMux
    port map (
            O => \N__49780\,
            I => \N__49716\
        );

    \I__11835\ : InMux
    port map (
            O => \N__49779\,
            I => \N__49716\
        );

    \I__11834\ : InMux
    port map (
            O => \N__49778\,
            I => \N__49716\
        );

    \I__11833\ : InMux
    port map (
            O => \N__49777\,
            I => \N__49716\
        );

    \I__11832\ : InMux
    port map (
            O => \N__49776\,
            I => \N__49711\
        );

    \I__11831\ : InMux
    port map (
            O => \N__49775\,
            I => \N__49711\
        );

    \I__11830\ : Span4Mux_v
    port map (
            O => \N__49772\,
            I => \N__49702\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__49767\,
            I => \N__49702\
        );

    \I__11828\ : InMux
    port map (
            O => \N__49766\,
            I => \N__49699\
        );

    \I__11827\ : InMux
    port map (
            O => \N__49765\,
            I => \N__49688\
        );

    \I__11826\ : InMux
    port map (
            O => \N__49764\,
            I => \N__49688\
        );

    \I__11825\ : InMux
    port map (
            O => \N__49763\,
            I => \N__49688\
        );

    \I__11824\ : InMux
    port map (
            O => \N__49762\,
            I => \N__49688\
        );

    \I__11823\ : InMux
    port map (
            O => \N__49761\,
            I => \N__49688\
        );

    \I__11822\ : LocalMux
    port map (
            O => \N__49758\,
            I => \N__49685\
        );

    \I__11821\ : InMux
    port map (
            O => \N__49757\,
            I => \N__49670\
        );

    \I__11820\ : InMux
    port map (
            O => \N__49756\,
            I => \N__49670\
        );

    \I__11819\ : InMux
    port map (
            O => \N__49755\,
            I => \N__49670\
        );

    \I__11818\ : InMux
    port map (
            O => \N__49754\,
            I => \N__49670\
        );

    \I__11817\ : InMux
    port map (
            O => \N__49753\,
            I => \N__49670\
        );

    \I__11816\ : InMux
    port map (
            O => \N__49752\,
            I => \N__49670\
        );

    \I__11815\ : InMux
    port map (
            O => \N__49751\,
            I => \N__49670\
        );

    \I__11814\ : InMux
    port map (
            O => \N__49750\,
            I => \N__49665\
        );

    \I__11813\ : InMux
    port map (
            O => \N__49749\,
            I => \N__49665\
        );

    \I__11812\ : InMux
    port map (
            O => \N__49748\,
            I => \N__49660\
        );

    \I__11811\ : InMux
    port map (
            O => \N__49747\,
            I => \N__49660\
        );

    \I__11810\ : InMux
    port map (
            O => \N__49746\,
            I => \N__49655\
        );

    \I__11809\ : InMux
    port map (
            O => \N__49745\,
            I => \N__49655\
        );

    \I__11808\ : InMux
    port map (
            O => \N__49744\,
            I => \N__49646\
        );

    \I__11807\ : InMux
    port map (
            O => \N__49743\,
            I => \N__49646\
        );

    \I__11806\ : InMux
    port map (
            O => \N__49742\,
            I => \N__49646\
        );

    \I__11805\ : InMux
    port map (
            O => \N__49741\,
            I => \N__49646\
        );

    \I__11804\ : InMux
    port map (
            O => \N__49740\,
            I => \N__49636\
        );

    \I__11803\ : InMux
    port map (
            O => \N__49739\,
            I => \N__49636\
        );

    \I__11802\ : InMux
    port map (
            O => \N__49738\,
            I => \N__49636\
        );

    \I__11801\ : InMux
    port map (
            O => \N__49737\,
            I => \N__49636\
        );

    \I__11800\ : InMux
    port map (
            O => \N__49736\,
            I => \N__49625\
        );

    \I__11799\ : InMux
    port map (
            O => \N__49735\,
            I => \N__49625\
        );

    \I__11798\ : InMux
    port map (
            O => \N__49734\,
            I => \N__49625\
        );

    \I__11797\ : InMux
    port map (
            O => \N__49733\,
            I => \N__49625\
        );

    \I__11796\ : InMux
    port map (
            O => \N__49732\,
            I => \N__49625\
        );

    \I__11795\ : LocalMux
    port map (
            O => \N__49729\,
            I => \N__49610\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__49716\,
            I => \N__49610\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__49711\,
            I => \N__49610\
        );

    \I__11792\ : InMux
    port map (
            O => \N__49710\,
            I => \N__49607\
        );

    \I__11791\ : InMux
    port map (
            O => \N__49709\,
            I => \N__49604\
        );

    \I__11790\ : InMux
    port map (
            O => \N__49708\,
            I => \N__49599\
        );

    \I__11789\ : InMux
    port map (
            O => \N__49707\,
            I => \N__49599\
        );

    \I__11788\ : Span4Mux_v
    port map (
            O => \N__49702\,
            I => \N__49596\
        );

    \I__11787\ : LocalMux
    port map (
            O => \N__49699\,
            I => \N__49591\
        );

    \I__11786\ : LocalMux
    port map (
            O => \N__49688\,
            I => \N__49591\
        );

    \I__11785\ : Span4Mux_v
    port map (
            O => \N__49685\,
            I => \N__49582\
        );

    \I__11784\ : LocalMux
    port map (
            O => \N__49670\,
            I => \N__49582\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__49665\,
            I => \N__49570\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__49660\,
            I => \N__49570\
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__49655\,
            I => \N__49570\
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__49646\,
            I => \N__49567\
        );

    \I__11779\ : CascadeMux
    port map (
            O => \N__49645\,
            I => \N__49562\
        );

    \I__11778\ : LocalMux
    port map (
            O => \N__49636\,
            I => \N__49556\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__49625\,
            I => \N__49556\
        );

    \I__11776\ : InMux
    port map (
            O => \N__49624\,
            I => \N__49539\
        );

    \I__11775\ : InMux
    port map (
            O => \N__49623\,
            I => \N__49539\
        );

    \I__11774\ : InMux
    port map (
            O => \N__49622\,
            I => \N__49539\
        );

    \I__11773\ : InMux
    port map (
            O => \N__49621\,
            I => \N__49539\
        );

    \I__11772\ : InMux
    port map (
            O => \N__49620\,
            I => \N__49539\
        );

    \I__11771\ : InMux
    port map (
            O => \N__49619\,
            I => \N__49539\
        );

    \I__11770\ : InMux
    port map (
            O => \N__49618\,
            I => \N__49539\
        );

    \I__11769\ : InMux
    port map (
            O => \N__49617\,
            I => \N__49539\
        );

    \I__11768\ : Span4Mux_v
    port map (
            O => \N__49610\,
            I => \N__49534\
        );

    \I__11767\ : LocalMux
    port map (
            O => \N__49607\,
            I => \N__49534\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__49604\,
            I => \N__49529\
        );

    \I__11765\ : LocalMux
    port map (
            O => \N__49599\,
            I => \N__49529\
        );

    \I__11764\ : Span4Mux_h
    port map (
            O => \N__49596\,
            I => \N__49526\
        );

    \I__11763\ : Span12Mux_s11_h
    port map (
            O => \N__49591\,
            I => \N__49523\
        );

    \I__11762\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49514\
        );

    \I__11761\ : InMux
    port map (
            O => \N__49589\,
            I => \N__49514\
        );

    \I__11760\ : InMux
    port map (
            O => \N__49588\,
            I => \N__49514\
        );

    \I__11759\ : InMux
    port map (
            O => \N__49587\,
            I => \N__49514\
        );

    \I__11758\ : Span4Mux_h
    port map (
            O => \N__49582\,
            I => \N__49511\
        );

    \I__11757\ : InMux
    port map (
            O => \N__49581\,
            I => \N__49508\
        );

    \I__11756\ : InMux
    port map (
            O => \N__49580\,
            I => \N__49499\
        );

    \I__11755\ : InMux
    port map (
            O => \N__49579\,
            I => \N__49499\
        );

    \I__11754\ : InMux
    port map (
            O => \N__49578\,
            I => \N__49499\
        );

    \I__11753\ : InMux
    port map (
            O => \N__49577\,
            I => \N__49499\
        );

    \I__11752\ : Span4Mux_h
    port map (
            O => \N__49570\,
            I => \N__49494\
        );

    \I__11751\ : Span4Mux_h
    port map (
            O => \N__49567\,
            I => \N__49494\
        );

    \I__11750\ : InMux
    port map (
            O => \N__49566\,
            I => \N__49485\
        );

    \I__11749\ : InMux
    port map (
            O => \N__49565\,
            I => \N__49485\
        );

    \I__11748\ : InMux
    port map (
            O => \N__49562\,
            I => \N__49485\
        );

    \I__11747\ : InMux
    port map (
            O => \N__49561\,
            I => \N__49485\
        );

    \I__11746\ : Span4Mux_v
    port map (
            O => \N__49556\,
            I => \N__49476\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__49539\,
            I => \N__49476\
        );

    \I__11744\ : Span4Mux_h
    port map (
            O => \N__49534\,
            I => \N__49476\
        );

    \I__11743\ : Span4Mux_v
    port map (
            O => \N__49529\,
            I => \N__49476\
        );

    \I__11742\ : Odrv4
    port map (
            O => \N__49526\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11741\ : Odrv12
    port map (
            O => \N__49523\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11740\ : LocalMux
    port map (
            O => \N__49514\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11739\ : Odrv4
    port map (
            O => \N__49511\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__49508\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11737\ : LocalMux
    port map (
            O => \N__49499\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11736\ : Odrv4
    port map (
            O => \N__49494\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__49485\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11734\ : Odrv4
    port map (
            O => \N__49476\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11733\ : CascadeMux
    port map (
            O => \N__49457\,
            I => \N__49451\
        );

    \I__11732\ : CascadeMux
    port map (
            O => \N__49456\,
            I => \N__49447\
        );

    \I__11731\ : CascadeMux
    port map (
            O => \N__49455\,
            I => \N__49444\
        );

    \I__11730\ : CascadeMux
    port map (
            O => \N__49454\,
            I => \N__49440\
        );

    \I__11729\ : InMux
    port map (
            O => \N__49451\,
            I => \N__49436\
        );

    \I__11728\ : CascadeMux
    port map (
            O => \N__49450\,
            I => \N__49424\
        );

    \I__11727\ : InMux
    port map (
            O => \N__49447\,
            I => \N__49420\
        );

    \I__11726\ : InMux
    port map (
            O => \N__49444\,
            I => \N__49417\
        );

    \I__11725\ : InMux
    port map (
            O => \N__49443\,
            I => \N__49414\
        );

    \I__11724\ : InMux
    port map (
            O => \N__49440\,
            I => \N__49409\
        );

    \I__11723\ : InMux
    port map (
            O => \N__49439\,
            I => \N__49409\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__49436\,
            I => \N__49406\
        );

    \I__11721\ : CascadeMux
    port map (
            O => \N__49435\,
            I => \N__49403\
        );

    \I__11720\ : CascadeMux
    port map (
            O => \N__49434\,
            I => \N__49397\
        );

    \I__11719\ : CascadeMux
    port map (
            O => \N__49433\,
            I => \N__49385\
        );

    \I__11718\ : CascadeMux
    port map (
            O => \N__49432\,
            I => \N__49382\
        );

    \I__11717\ : CascadeMux
    port map (
            O => \N__49431\,
            I => \N__49374\
        );

    \I__11716\ : CascadeMux
    port map (
            O => \N__49430\,
            I => \N__49371\
        );

    \I__11715\ : CascadeMux
    port map (
            O => \N__49429\,
            I => \N__49366\
        );

    \I__11714\ : CascadeMux
    port map (
            O => \N__49428\,
            I => \N__49363\
        );

    \I__11713\ : InMux
    port map (
            O => \N__49427\,
            I => \N__49342\
        );

    \I__11712\ : InMux
    port map (
            O => \N__49424\,
            I => \N__49342\
        );

    \I__11711\ : InMux
    port map (
            O => \N__49423\,
            I => \N__49342\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__49420\,
            I => \N__49337\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__49417\,
            I => \N__49337\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__49414\,
            I => \N__49332\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__49409\,
            I => \N__49332\
        );

    \I__11706\ : Span4Mux_h
    port map (
            O => \N__49406\,
            I => \N__49329\
        );

    \I__11705\ : InMux
    port map (
            O => \N__49403\,
            I => \N__49318\
        );

    \I__11704\ : InMux
    port map (
            O => \N__49402\,
            I => \N__49318\
        );

    \I__11703\ : InMux
    port map (
            O => \N__49401\,
            I => \N__49318\
        );

    \I__11702\ : InMux
    port map (
            O => \N__49400\,
            I => \N__49318\
        );

    \I__11701\ : InMux
    port map (
            O => \N__49397\,
            I => \N__49318\
        );

    \I__11700\ : CascadeMux
    port map (
            O => \N__49396\,
            I => \N__49315\
        );

    \I__11699\ : CascadeMux
    port map (
            O => \N__49395\,
            I => \N__49312\
        );

    \I__11698\ : CascadeMux
    port map (
            O => \N__49394\,
            I => \N__49305\
        );

    \I__11697\ : CascadeMux
    port map (
            O => \N__49393\,
            I => \N__49302\
        );

    \I__11696\ : CascadeMux
    port map (
            O => \N__49392\,
            I => \N__49299\
        );

    \I__11695\ : CascadeMux
    port map (
            O => \N__49391\,
            I => \N__49296\
        );

    \I__11694\ : CascadeMux
    port map (
            O => \N__49390\,
            I => \N__49293\
        );

    \I__11693\ : CascadeMux
    port map (
            O => \N__49389\,
            I => \N__49289\
        );

    \I__11692\ : CascadeMux
    port map (
            O => \N__49388\,
            I => \N__49286\
        );

    \I__11691\ : InMux
    port map (
            O => \N__49385\,
            I => \N__49267\
        );

    \I__11690\ : InMux
    port map (
            O => \N__49382\,
            I => \N__49267\
        );

    \I__11689\ : CascadeMux
    port map (
            O => \N__49381\,
            I => \N__49263\
        );

    \I__11688\ : CascadeMux
    port map (
            O => \N__49380\,
            I => \N__49260\
        );

    \I__11687\ : CascadeMux
    port map (
            O => \N__49379\,
            I => \N__49257\
        );

    \I__11686\ : CascadeMux
    port map (
            O => \N__49378\,
            I => \N__49251\
        );

    \I__11685\ : InMux
    port map (
            O => \N__49377\,
            I => \N__49243\
        );

    \I__11684\ : InMux
    port map (
            O => \N__49374\,
            I => \N__49243\
        );

    \I__11683\ : InMux
    port map (
            O => \N__49371\,
            I => \N__49236\
        );

    \I__11682\ : InMux
    port map (
            O => \N__49370\,
            I => \N__49236\
        );

    \I__11681\ : InMux
    port map (
            O => \N__49369\,
            I => \N__49236\
        );

    \I__11680\ : InMux
    port map (
            O => \N__49366\,
            I => \N__49231\
        );

    \I__11679\ : InMux
    port map (
            O => \N__49363\,
            I => \N__49231\
        );

    \I__11678\ : CascadeMux
    port map (
            O => \N__49362\,
            I => \N__49228\
        );

    \I__11677\ : CascadeMux
    port map (
            O => \N__49361\,
            I => \N__49225\
        );

    \I__11676\ : CascadeMux
    port map (
            O => \N__49360\,
            I => \N__49221\
        );

    \I__11675\ : CascadeMux
    port map (
            O => \N__49359\,
            I => \N__49217\
        );

    \I__11674\ : CascadeMux
    port map (
            O => \N__49358\,
            I => \N__49213\
        );

    \I__11673\ : CascadeMux
    port map (
            O => \N__49357\,
            I => \N__49209\
        );

    \I__11672\ : CascadeMux
    port map (
            O => \N__49356\,
            I => \N__49205\
        );

    \I__11671\ : CascadeMux
    port map (
            O => \N__49355\,
            I => \N__49192\
        );

    \I__11670\ : CascadeMux
    port map (
            O => \N__49354\,
            I => \N__49188\
        );

    \I__11669\ : CascadeMux
    port map (
            O => \N__49353\,
            I => \N__49184\
        );

    \I__11668\ : CascadeMux
    port map (
            O => \N__49352\,
            I => \N__49180\
        );

    \I__11667\ : CascadeMux
    port map (
            O => \N__49351\,
            I => \N__49175\
        );

    \I__11666\ : CascadeMux
    port map (
            O => \N__49350\,
            I => \N__49171\
        );

    \I__11665\ : CascadeMux
    port map (
            O => \N__49349\,
            I => \N__49167\
        );

    \I__11664\ : LocalMux
    port map (
            O => \N__49342\,
            I => \N__49164\
        );

    \I__11663\ : Span4Mux_v
    port map (
            O => \N__49337\,
            I => \N__49159\
        );

    \I__11662\ : Span4Mux_v
    port map (
            O => \N__49332\,
            I => \N__49159\
        );

    \I__11661\ : Span4Mux_h
    port map (
            O => \N__49329\,
            I => \N__49154\
        );

    \I__11660\ : LocalMux
    port map (
            O => \N__49318\,
            I => \N__49154\
        );

    \I__11659\ : InMux
    port map (
            O => \N__49315\,
            I => \N__49137\
        );

    \I__11658\ : InMux
    port map (
            O => \N__49312\,
            I => \N__49137\
        );

    \I__11657\ : InMux
    port map (
            O => \N__49311\,
            I => \N__49137\
        );

    \I__11656\ : InMux
    port map (
            O => \N__49310\,
            I => \N__49137\
        );

    \I__11655\ : InMux
    port map (
            O => \N__49309\,
            I => \N__49137\
        );

    \I__11654\ : InMux
    port map (
            O => \N__49308\,
            I => \N__49137\
        );

    \I__11653\ : InMux
    port map (
            O => \N__49305\,
            I => \N__49137\
        );

    \I__11652\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49137\
        );

    \I__11651\ : InMux
    port map (
            O => \N__49299\,
            I => \N__49128\
        );

    \I__11650\ : InMux
    port map (
            O => \N__49296\,
            I => \N__49128\
        );

    \I__11649\ : InMux
    port map (
            O => \N__49293\,
            I => \N__49128\
        );

    \I__11648\ : InMux
    port map (
            O => \N__49292\,
            I => \N__49128\
        );

    \I__11647\ : InMux
    port map (
            O => \N__49289\,
            I => \N__49123\
        );

    \I__11646\ : InMux
    port map (
            O => \N__49286\,
            I => \N__49123\
        );

    \I__11645\ : CascadeMux
    port map (
            O => \N__49285\,
            I => \N__49120\
        );

    \I__11644\ : CascadeMux
    port map (
            O => \N__49284\,
            I => \N__49117\
        );

    \I__11643\ : CascadeMux
    port map (
            O => \N__49283\,
            I => \N__49114\
        );

    \I__11642\ : CascadeMux
    port map (
            O => \N__49282\,
            I => \N__49111\
        );

    \I__11641\ : CascadeMux
    port map (
            O => \N__49281\,
            I => \N__49107\
        );

    \I__11640\ : CascadeMux
    port map (
            O => \N__49280\,
            I => \N__49100\
        );

    \I__11639\ : CascadeMux
    port map (
            O => \N__49279\,
            I => \N__49096\
        );

    \I__11638\ : CascadeMux
    port map (
            O => \N__49278\,
            I => \N__49092\
        );

    \I__11637\ : CascadeMux
    port map (
            O => \N__49277\,
            I => \N__49088\
        );

    \I__11636\ : CascadeMux
    port map (
            O => \N__49276\,
            I => \N__49084\
        );

    \I__11635\ : CascadeMux
    port map (
            O => \N__49275\,
            I => \N__49081\
        );

    \I__11634\ : CascadeMux
    port map (
            O => \N__49274\,
            I => \N__49077\
        );

    \I__11633\ : CascadeMux
    port map (
            O => \N__49273\,
            I => \N__49073\
        );

    \I__11632\ : CascadeMux
    port map (
            O => \N__49272\,
            I => \N__49069\
        );

    \I__11631\ : LocalMux
    port map (
            O => \N__49267\,
            I => \N__49065\
        );

    \I__11630\ : InMux
    port map (
            O => \N__49266\,
            I => \N__49060\
        );

    \I__11629\ : InMux
    port map (
            O => \N__49263\,
            I => \N__49060\
        );

    \I__11628\ : InMux
    port map (
            O => \N__49260\,
            I => \N__49055\
        );

    \I__11627\ : InMux
    port map (
            O => \N__49257\,
            I => \N__49055\
        );

    \I__11626\ : InMux
    port map (
            O => \N__49256\,
            I => \N__49040\
        );

    \I__11625\ : InMux
    port map (
            O => \N__49255\,
            I => \N__49040\
        );

    \I__11624\ : InMux
    port map (
            O => \N__49254\,
            I => \N__49040\
        );

    \I__11623\ : InMux
    port map (
            O => \N__49251\,
            I => \N__49040\
        );

    \I__11622\ : InMux
    port map (
            O => \N__49250\,
            I => \N__49040\
        );

    \I__11621\ : InMux
    port map (
            O => \N__49249\,
            I => \N__49040\
        );

    \I__11620\ : InMux
    port map (
            O => \N__49248\,
            I => \N__49040\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__49243\,
            I => \N__49035\
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__49236\,
            I => \N__49035\
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__49231\,
            I => \N__49032\
        );

    \I__11616\ : InMux
    port map (
            O => \N__49228\,
            I => \N__49021\
        );

    \I__11615\ : InMux
    port map (
            O => \N__49225\,
            I => \N__49021\
        );

    \I__11614\ : InMux
    port map (
            O => \N__49224\,
            I => \N__49021\
        );

    \I__11613\ : InMux
    port map (
            O => \N__49221\,
            I => \N__49021\
        );

    \I__11612\ : InMux
    port map (
            O => \N__49220\,
            I => \N__49021\
        );

    \I__11611\ : InMux
    port map (
            O => \N__49217\,
            I => \N__49004\
        );

    \I__11610\ : InMux
    port map (
            O => \N__49216\,
            I => \N__49004\
        );

    \I__11609\ : InMux
    port map (
            O => \N__49213\,
            I => \N__49004\
        );

    \I__11608\ : InMux
    port map (
            O => \N__49212\,
            I => \N__49004\
        );

    \I__11607\ : InMux
    port map (
            O => \N__49209\,
            I => \N__49004\
        );

    \I__11606\ : InMux
    port map (
            O => \N__49208\,
            I => \N__49004\
        );

    \I__11605\ : InMux
    port map (
            O => \N__49205\,
            I => \N__49004\
        );

    \I__11604\ : InMux
    port map (
            O => \N__49204\,
            I => \N__49004\
        );

    \I__11603\ : CascadeMux
    port map (
            O => \N__49203\,
            I => \N__49001\
        );

    \I__11602\ : CascadeMux
    port map (
            O => \N__49202\,
            I => \N__48998\
        );

    \I__11601\ : CascadeMux
    port map (
            O => \N__49201\,
            I => \N__48995\
        );

    \I__11600\ : CascadeMux
    port map (
            O => \N__49200\,
            I => \N__48991\
        );

    \I__11599\ : CascadeMux
    port map (
            O => \N__49199\,
            I => \N__48988\
        );

    \I__11598\ : CascadeMux
    port map (
            O => \N__49198\,
            I => \N__48985\
        );

    \I__11597\ : CascadeMux
    port map (
            O => \N__49197\,
            I => \N__48980\
        );

    \I__11596\ : CascadeMux
    port map (
            O => \N__49196\,
            I => \N__48976\
        );

    \I__11595\ : CascadeMux
    port map (
            O => \N__49195\,
            I => \N__48972\
        );

    \I__11594\ : InMux
    port map (
            O => \N__49192\,
            I => \N__48955\
        );

    \I__11593\ : InMux
    port map (
            O => \N__49191\,
            I => \N__48955\
        );

    \I__11592\ : InMux
    port map (
            O => \N__49188\,
            I => \N__48955\
        );

    \I__11591\ : InMux
    port map (
            O => \N__49187\,
            I => \N__48955\
        );

    \I__11590\ : InMux
    port map (
            O => \N__49184\,
            I => \N__48955\
        );

    \I__11589\ : InMux
    port map (
            O => \N__49183\,
            I => \N__48955\
        );

    \I__11588\ : InMux
    port map (
            O => \N__49180\,
            I => \N__48955\
        );

    \I__11587\ : InMux
    port map (
            O => \N__49179\,
            I => \N__48955\
        );

    \I__11586\ : InMux
    port map (
            O => \N__49178\,
            I => \N__48942\
        );

    \I__11585\ : InMux
    port map (
            O => \N__49175\,
            I => \N__48942\
        );

    \I__11584\ : InMux
    port map (
            O => \N__49174\,
            I => \N__48942\
        );

    \I__11583\ : InMux
    port map (
            O => \N__49171\,
            I => \N__48942\
        );

    \I__11582\ : InMux
    port map (
            O => \N__49170\,
            I => \N__48942\
        );

    \I__11581\ : InMux
    port map (
            O => \N__49167\,
            I => \N__48942\
        );

    \I__11580\ : Span4Mux_h
    port map (
            O => \N__49164\,
            I => \N__48939\
        );

    \I__11579\ : Sp12to4
    port map (
            O => \N__49159\,
            I => \N__48936\
        );

    \I__11578\ : Span4Mux_h
    port map (
            O => \N__49154\,
            I => \N__48931\
        );

    \I__11577\ : LocalMux
    port map (
            O => \N__49137\,
            I => \N__48931\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__49128\,
            I => \N__48926\
        );

    \I__11575\ : LocalMux
    port map (
            O => \N__49123\,
            I => \N__48926\
        );

    \I__11574\ : InMux
    port map (
            O => \N__49120\,
            I => \N__48917\
        );

    \I__11573\ : InMux
    port map (
            O => \N__49117\,
            I => \N__48917\
        );

    \I__11572\ : InMux
    port map (
            O => \N__49114\,
            I => \N__48917\
        );

    \I__11571\ : InMux
    port map (
            O => \N__49111\,
            I => \N__48917\
        );

    \I__11570\ : InMux
    port map (
            O => \N__49110\,
            I => \N__48912\
        );

    \I__11569\ : InMux
    port map (
            O => \N__49107\,
            I => \N__48912\
        );

    \I__11568\ : InMux
    port map (
            O => \N__49106\,
            I => \N__48903\
        );

    \I__11567\ : InMux
    port map (
            O => \N__49105\,
            I => \N__48903\
        );

    \I__11566\ : InMux
    port map (
            O => \N__49104\,
            I => \N__48903\
        );

    \I__11565\ : InMux
    port map (
            O => \N__49103\,
            I => \N__48903\
        );

    \I__11564\ : InMux
    port map (
            O => \N__49100\,
            I => \N__48900\
        );

    \I__11563\ : InMux
    port map (
            O => \N__49099\,
            I => \N__48883\
        );

    \I__11562\ : InMux
    port map (
            O => \N__49096\,
            I => \N__48883\
        );

    \I__11561\ : InMux
    port map (
            O => \N__49095\,
            I => \N__48883\
        );

    \I__11560\ : InMux
    port map (
            O => \N__49092\,
            I => \N__48883\
        );

    \I__11559\ : InMux
    port map (
            O => \N__49091\,
            I => \N__48883\
        );

    \I__11558\ : InMux
    port map (
            O => \N__49088\,
            I => \N__48883\
        );

    \I__11557\ : InMux
    port map (
            O => \N__49087\,
            I => \N__48883\
        );

    \I__11556\ : InMux
    port map (
            O => \N__49084\,
            I => \N__48883\
        );

    \I__11555\ : InMux
    port map (
            O => \N__49081\,
            I => \N__48866\
        );

    \I__11554\ : InMux
    port map (
            O => \N__49080\,
            I => \N__48866\
        );

    \I__11553\ : InMux
    port map (
            O => \N__49077\,
            I => \N__48866\
        );

    \I__11552\ : InMux
    port map (
            O => \N__49076\,
            I => \N__48866\
        );

    \I__11551\ : InMux
    port map (
            O => \N__49073\,
            I => \N__48866\
        );

    \I__11550\ : InMux
    port map (
            O => \N__49072\,
            I => \N__48866\
        );

    \I__11549\ : InMux
    port map (
            O => \N__49069\,
            I => \N__48866\
        );

    \I__11548\ : InMux
    port map (
            O => \N__49068\,
            I => \N__48866\
        );

    \I__11547\ : Span4Mux_v
    port map (
            O => \N__49065\,
            I => \N__48849\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__49060\,
            I => \N__48849\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__49055\,
            I => \N__48849\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__49040\,
            I => \N__48849\
        );

    \I__11543\ : Span4Mux_h
    port map (
            O => \N__49035\,
            I => \N__48849\
        );

    \I__11542\ : Span4Mux_h
    port map (
            O => \N__49032\,
            I => \N__48849\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__49021\,
            I => \N__48849\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__49004\,
            I => \N__48849\
        );

    \I__11539\ : InMux
    port map (
            O => \N__49001\,
            I => \N__48840\
        );

    \I__11538\ : InMux
    port map (
            O => \N__48998\,
            I => \N__48840\
        );

    \I__11537\ : InMux
    port map (
            O => \N__48995\,
            I => \N__48840\
        );

    \I__11536\ : InMux
    port map (
            O => \N__48994\,
            I => \N__48840\
        );

    \I__11535\ : InMux
    port map (
            O => \N__48991\,
            I => \N__48831\
        );

    \I__11534\ : InMux
    port map (
            O => \N__48988\,
            I => \N__48831\
        );

    \I__11533\ : InMux
    port map (
            O => \N__48985\,
            I => \N__48831\
        );

    \I__11532\ : InMux
    port map (
            O => \N__48984\,
            I => \N__48831\
        );

    \I__11531\ : InMux
    port map (
            O => \N__48983\,
            I => \N__48818\
        );

    \I__11530\ : InMux
    port map (
            O => \N__48980\,
            I => \N__48818\
        );

    \I__11529\ : InMux
    port map (
            O => \N__48979\,
            I => \N__48818\
        );

    \I__11528\ : InMux
    port map (
            O => \N__48976\,
            I => \N__48818\
        );

    \I__11527\ : InMux
    port map (
            O => \N__48975\,
            I => \N__48818\
        );

    \I__11526\ : InMux
    port map (
            O => \N__48972\,
            I => \N__48818\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__48955\,
            I => \N__48813\
        );

    \I__11524\ : LocalMux
    port map (
            O => \N__48942\,
            I => \N__48813\
        );

    \I__11523\ : Odrv4
    port map (
            O => \N__48939\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11522\ : Odrv12
    port map (
            O => \N__48936\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11521\ : Odrv4
    port map (
            O => \N__48931\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11520\ : Odrv4
    port map (
            O => \N__48926\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__48917\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__48912\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__48903\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__48900\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__48883\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11514\ : LocalMux
    port map (
            O => \N__48866\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11513\ : Odrv4
    port map (
            O => \N__48849\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11512\ : LocalMux
    port map (
            O => \N__48840\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11511\ : LocalMux
    port map (
            O => \N__48831\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__48818\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11509\ : Odrv4
    port map (
            O => \N__48813\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11508\ : InMux
    port map (
            O => \N__48782\,
            I => \N__48779\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__48779\,
            I => \N__48776\
        );

    \I__11506\ : Span4Mux_h
    port map (
            O => \N__48776\,
            I => \N__48773\
        );

    \I__11505\ : Odrv4
    port map (
            O => \N__48773\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__11504\ : InMux
    port map (
            O => \N__48770\,
            I => \N__48765\
        );

    \I__11503\ : InMux
    port map (
            O => \N__48769\,
            I => \N__48760\
        );

    \I__11502\ : InMux
    port map (
            O => \N__48768\,
            I => \N__48760\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__48765\,
            I => \N__48755\
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__48760\,
            I => \N__48755\
        );

    \I__11499\ : Span4Mux_h
    port map (
            O => \N__48755\,
            I => \N__48751\
        );

    \I__11498\ : InMux
    port map (
            O => \N__48754\,
            I => \N__48748\
        );

    \I__11497\ : Odrv4
    port map (
            O => \N__48751\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__48748\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__11495\ : InMux
    port map (
            O => \N__48743\,
            I => \N__48734\
        );

    \I__11494\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48734\
        );

    \I__11493\ : InMux
    port map (
            O => \N__48741\,
            I => \N__48734\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__48734\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__11491\ : InMux
    port map (
            O => \N__48731\,
            I => \N__48728\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__48728\,
            I => \N__48725\
        );

    \I__11489\ : Odrv12
    port map (
            O => \N__48725\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__11488\ : InMux
    port map (
            O => \N__48722\,
            I => \N__48718\
        );

    \I__11487\ : InMux
    port map (
            O => \N__48721\,
            I => \N__48715\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__48718\,
            I => \N__48712\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__48715\,
            I => \N__48709\
        );

    \I__11484\ : Span4Mux_h
    port map (
            O => \N__48712\,
            I => \N__48706\
        );

    \I__11483\ : Span4Mux_h
    port map (
            O => \N__48709\,
            I => \N__48702\
        );

    \I__11482\ : Span4Mux_v
    port map (
            O => \N__48706\,
            I => \N__48699\
        );

    \I__11481\ : InMux
    port map (
            O => \N__48705\,
            I => \N__48696\
        );

    \I__11480\ : Odrv4
    port map (
            O => \N__48702\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__11479\ : Odrv4
    port map (
            O => \N__48699\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__48696\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__11477\ : InMux
    port map (
            O => \N__48689\,
            I => \N__48680\
        );

    \I__11476\ : InMux
    port map (
            O => \N__48688\,
            I => \N__48680\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48687\,
            I => \N__48677\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48686\,
            I => \N__48662\
        );

    \I__11473\ : CascadeMux
    port map (
            O => \N__48685\,
            I => \N__48659\
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__48680\,
            I => \N__48653\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__48677\,
            I => \N__48653\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48676\,
            I => \N__48640\
        );

    \I__11469\ : InMux
    port map (
            O => \N__48675\,
            I => \N__48640\
        );

    \I__11468\ : InMux
    port map (
            O => \N__48674\,
            I => \N__48640\
        );

    \I__11467\ : InMux
    port map (
            O => \N__48673\,
            I => \N__48640\
        );

    \I__11466\ : InMux
    port map (
            O => \N__48672\,
            I => \N__48640\
        );

    \I__11465\ : InMux
    port map (
            O => \N__48671\,
            I => \N__48640\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48670\,
            I => \N__48635\
        );

    \I__11463\ : InMux
    port map (
            O => \N__48669\,
            I => \N__48635\
        );

    \I__11462\ : InMux
    port map (
            O => \N__48668\,
            I => \N__48630\
        );

    \I__11461\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48630\
        );

    \I__11460\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48625\
        );

    \I__11459\ : InMux
    port map (
            O => \N__48665\,
            I => \N__48625\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__48662\,
            I => \N__48622\
        );

    \I__11457\ : InMux
    port map (
            O => \N__48659\,
            I => \N__48617\
        );

    \I__11456\ : InMux
    port map (
            O => \N__48658\,
            I => \N__48617\
        );

    \I__11455\ : Span4Mux_v
    port map (
            O => \N__48653\,
            I => \N__48614\
        );

    \I__11454\ : LocalMux
    port map (
            O => \N__48640\,
            I => \N__48609\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__48635\,
            I => \N__48609\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__48630\,
            I => \N__48598\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__48625\,
            I => \N__48598\
        );

    \I__11450\ : Span4Mux_h
    port map (
            O => \N__48622\,
            I => \N__48595\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__48617\,
            I => \N__48588\
        );

    \I__11448\ : Span4Mux_h
    port map (
            O => \N__48614\,
            I => \N__48588\
        );

    \I__11447\ : Span4Mux_v
    port map (
            O => \N__48609\,
            I => \N__48588\
        );

    \I__11446\ : InMux
    port map (
            O => \N__48608\,
            I => \N__48579\
        );

    \I__11445\ : InMux
    port map (
            O => \N__48607\,
            I => \N__48579\
        );

    \I__11444\ : InMux
    port map (
            O => \N__48606\,
            I => \N__48579\
        );

    \I__11443\ : InMux
    port map (
            O => \N__48605\,
            I => \N__48579\
        );

    \I__11442\ : InMux
    port map (
            O => \N__48604\,
            I => \N__48576\
        );

    \I__11441\ : InMux
    port map (
            O => \N__48603\,
            I => \N__48572\
        );

    \I__11440\ : Span4Mux_v
    port map (
            O => \N__48598\,
            I => \N__48569\
        );

    \I__11439\ : Span4Mux_v
    port map (
            O => \N__48595\,
            I => \N__48566\
        );

    \I__11438\ : Sp12to4
    port map (
            O => \N__48588\,
            I => \N__48559\
        );

    \I__11437\ : LocalMux
    port map (
            O => \N__48579\,
            I => \N__48559\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__48576\,
            I => \N__48559\
        );

    \I__11435\ : InMux
    port map (
            O => \N__48575\,
            I => \N__48556\
        );

    \I__11434\ : LocalMux
    port map (
            O => \N__48572\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__11433\ : Odrv4
    port map (
            O => \N__48569\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__11432\ : Odrv4
    port map (
            O => \N__48566\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__11431\ : Odrv12
    port map (
            O => \N__48559\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__11430\ : LocalMux
    port map (
            O => \N__48556\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__11429\ : CascadeMux
    port map (
            O => \N__48545\,
            I => \N__48541\
        );

    \I__11428\ : InMux
    port map (
            O => \N__48544\,
            I => \N__48538\
        );

    \I__11427\ : InMux
    port map (
            O => \N__48541\,
            I => \N__48535\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__48538\,
            I => \N__48532\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__48535\,
            I => \N__48528\
        );

    \I__11424\ : Span12Mux_s10_h
    port map (
            O => \N__48532\,
            I => \N__48525\
        );

    \I__11423\ : InMux
    port map (
            O => \N__48531\,
            I => \N__48522\
        );

    \I__11422\ : Span4Mux_v
    port map (
            O => \N__48528\,
            I => \N__48519\
        );

    \I__11421\ : Odrv12
    port map (
            O => \N__48525\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__48522\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__11419\ : Odrv4
    port map (
            O => \N__48519\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__11418\ : InMux
    port map (
            O => \N__48512\,
            I => \N__48509\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__48509\,
            I => \N__48505\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48508\,
            I => \N__48502\
        );

    \I__11415\ : Span4Mux_h
    port map (
            O => \N__48505\,
            I => \N__48497\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__48502\,
            I => \N__48497\
        );

    \I__11413\ : Span4Mux_v
    port map (
            O => \N__48497\,
            I => \N__48492\
        );

    \I__11412\ : InMux
    port map (
            O => \N__48496\,
            I => \N__48487\
        );

    \I__11411\ : InMux
    port map (
            O => \N__48495\,
            I => \N__48487\
        );

    \I__11410\ : Odrv4
    port map (
            O => \N__48492\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__48487\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__11408\ : ClkMux
    port map (
            O => \N__48482\,
            I => \N__48020\
        );

    \I__11407\ : ClkMux
    port map (
            O => \N__48481\,
            I => \N__48020\
        );

    \I__11406\ : ClkMux
    port map (
            O => \N__48480\,
            I => \N__48020\
        );

    \I__11405\ : ClkMux
    port map (
            O => \N__48479\,
            I => \N__48020\
        );

    \I__11404\ : ClkMux
    port map (
            O => \N__48478\,
            I => \N__48020\
        );

    \I__11403\ : ClkMux
    port map (
            O => \N__48477\,
            I => \N__48020\
        );

    \I__11402\ : ClkMux
    port map (
            O => \N__48476\,
            I => \N__48020\
        );

    \I__11401\ : ClkMux
    port map (
            O => \N__48475\,
            I => \N__48020\
        );

    \I__11400\ : ClkMux
    port map (
            O => \N__48474\,
            I => \N__48020\
        );

    \I__11399\ : ClkMux
    port map (
            O => \N__48473\,
            I => \N__48020\
        );

    \I__11398\ : ClkMux
    port map (
            O => \N__48472\,
            I => \N__48020\
        );

    \I__11397\ : ClkMux
    port map (
            O => \N__48471\,
            I => \N__48020\
        );

    \I__11396\ : ClkMux
    port map (
            O => \N__48470\,
            I => \N__48020\
        );

    \I__11395\ : ClkMux
    port map (
            O => \N__48469\,
            I => \N__48020\
        );

    \I__11394\ : ClkMux
    port map (
            O => \N__48468\,
            I => \N__48020\
        );

    \I__11393\ : ClkMux
    port map (
            O => \N__48467\,
            I => \N__48020\
        );

    \I__11392\ : ClkMux
    port map (
            O => \N__48466\,
            I => \N__48020\
        );

    \I__11391\ : ClkMux
    port map (
            O => \N__48465\,
            I => \N__48020\
        );

    \I__11390\ : ClkMux
    port map (
            O => \N__48464\,
            I => \N__48020\
        );

    \I__11389\ : ClkMux
    port map (
            O => \N__48463\,
            I => \N__48020\
        );

    \I__11388\ : ClkMux
    port map (
            O => \N__48462\,
            I => \N__48020\
        );

    \I__11387\ : ClkMux
    port map (
            O => \N__48461\,
            I => \N__48020\
        );

    \I__11386\ : ClkMux
    port map (
            O => \N__48460\,
            I => \N__48020\
        );

    \I__11385\ : ClkMux
    port map (
            O => \N__48459\,
            I => \N__48020\
        );

    \I__11384\ : ClkMux
    port map (
            O => \N__48458\,
            I => \N__48020\
        );

    \I__11383\ : ClkMux
    port map (
            O => \N__48457\,
            I => \N__48020\
        );

    \I__11382\ : ClkMux
    port map (
            O => \N__48456\,
            I => \N__48020\
        );

    \I__11381\ : ClkMux
    port map (
            O => \N__48455\,
            I => \N__48020\
        );

    \I__11380\ : ClkMux
    port map (
            O => \N__48454\,
            I => \N__48020\
        );

    \I__11379\ : ClkMux
    port map (
            O => \N__48453\,
            I => \N__48020\
        );

    \I__11378\ : ClkMux
    port map (
            O => \N__48452\,
            I => \N__48020\
        );

    \I__11377\ : ClkMux
    port map (
            O => \N__48451\,
            I => \N__48020\
        );

    \I__11376\ : ClkMux
    port map (
            O => \N__48450\,
            I => \N__48020\
        );

    \I__11375\ : ClkMux
    port map (
            O => \N__48449\,
            I => \N__48020\
        );

    \I__11374\ : ClkMux
    port map (
            O => \N__48448\,
            I => \N__48020\
        );

    \I__11373\ : ClkMux
    port map (
            O => \N__48447\,
            I => \N__48020\
        );

    \I__11372\ : ClkMux
    port map (
            O => \N__48446\,
            I => \N__48020\
        );

    \I__11371\ : ClkMux
    port map (
            O => \N__48445\,
            I => \N__48020\
        );

    \I__11370\ : ClkMux
    port map (
            O => \N__48444\,
            I => \N__48020\
        );

    \I__11369\ : ClkMux
    port map (
            O => \N__48443\,
            I => \N__48020\
        );

    \I__11368\ : ClkMux
    port map (
            O => \N__48442\,
            I => \N__48020\
        );

    \I__11367\ : ClkMux
    port map (
            O => \N__48441\,
            I => \N__48020\
        );

    \I__11366\ : ClkMux
    port map (
            O => \N__48440\,
            I => \N__48020\
        );

    \I__11365\ : ClkMux
    port map (
            O => \N__48439\,
            I => \N__48020\
        );

    \I__11364\ : ClkMux
    port map (
            O => \N__48438\,
            I => \N__48020\
        );

    \I__11363\ : ClkMux
    port map (
            O => \N__48437\,
            I => \N__48020\
        );

    \I__11362\ : ClkMux
    port map (
            O => \N__48436\,
            I => \N__48020\
        );

    \I__11361\ : ClkMux
    port map (
            O => \N__48435\,
            I => \N__48020\
        );

    \I__11360\ : ClkMux
    port map (
            O => \N__48434\,
            I => \N__48020\
        );

    \I__11359\ : ClkMux
    port map (
            O => \N__48433\,
            I => \N__48020\
        );

    \I__11358\ : ClkMux
    port map (
            O => \N__48432\,
            I => \N__48020\
        );

    \I__11357\ : ClkMux
    port map (
            O => \N__48431\,
            I => \N__48020\
        );

    \I__11356\ : ClkMux
    port map (
            O => \N__48430\,
            I => \N__48020\
        );

    \I__11355\ : ClkMux
    port map (
            O => \N__48429\,
            I => \N__48020\
        );

    \I__11354\ : ClkMux
    port map (
            O => \N__48428\,
            I => \N__48020\
        );

    \I__11353\ : ClkMux
    port map (
            O => \N__48427\,
            I => \N__48020\
        );

    \I__11352\ : ClkMux
    port map (
            O => \N__48426\,
            I => \N__48020\
        );

    \I__11351\ : ClkMux
    port map (
            O => \N__48425\,
            I => \N__48020\
        );

    \I__11350\ : ClkMux
    port map (
            O => \N__48424\,
            I => \N__48020\
        );

    \I__11349\ : ClkMux
    port map (
            O => \N__48423\,
            I => \N__48020\
        );

    \I__11348\ : ClkMux
    port map (
            O => \N__48422\,
            I => \N__48020\
        );

    \I__11347\ : ClkMux
    port map (
            O => \N__48421\,
            I => \N__48020\
        );

    \I__11346\ : ClkMux
    port map (
            O => \N__48420\,
            I => \N__48020\
        );

    \I__11345\ : ClkMux
    port map (
            O => \N__48419\,
            I => \N__48020\
        );

    \I__11344\ : ClkMux
    port map (
            O => \N__48418\,
            I => \N__48020\
        );

    \I__11343\ : ClkMux
    port map (
            O => \N__48417\,
            I => \N__48020\
        );

    \I__11342\ : ClkMux
    port map (
            O => \N__48416\,
            I => \N__48020\
        );

    \I__11341\ : ClkMux
    port map (
            O => \N__48415\,
            I => \N__48020\
        );

    \I__11340\ : ClkMux
    port map (
            O => \N__48414\,
            I => \N__48020\
        );

    \I__11339\ : ClkMux
    port map (
            O => \N__48413\,
            I => \N__48020\
        );

    \I__11338\ : ClkMux
    port map (
            O => \N__48412\,
            I => \N__48020\
        );

    \I__11337\ : ClkMux
    port map (
            O => \N__48411\,
            I => \N__48020\
        );

    \I__11336\ : ClkMux
    port map (
            O => \N__48410\,
            I => \N__48020\
        );

    \I__11335\ : ClkMux
    port map (
            O => \N__48409\,
            I => \N__48020\
        );

    \I__11334\ : ClkMux
    port map (
            O => \N__48408\,
            I => \N__48020\
        );

    \I__11333\ : ClkMux
    port map (
            O => \N__48407\,
            I => \N__48020\
        );

    \I__11332\ : ClkMux
    port map (
            O => \N__48406\,
            I => \N__48020\
        );

    \I__11331\ : ClkMux
    port map (
            O => \N__48405\,
            I => \N__48020\
        );

    \I__11330\ : ClkMux
    port map (
            O => \N__48404\,
            I => \N__48020\
        );

    \I__11329\ : ClkMux
    port map (
            O => \N__48403\,
            I => \N__48020\
        );

    \I__11328\ : ClkMux
    port map (
            O => \N__48402\,
            I => \N__48020\
        );

    \I__11327\ : ClkMux
    port map (
            O => \N__48401\,
            I => \N__48020\
        );

    \I__11326\ : ClkMux
    port map (
            O => \N__48400\,
            I => \N__48020\
        );

    \I__11325\ : ClkMux
    port map (
            O => \N__48399\,
            I => \N__48020\
        );

    \I__11324\ : ClkMux
    port map (
            O => \N__48398\,
            I => \N__48020\
        );

    \I__11323\ : ClkMux
    port map (
            O => \N__48397\,
            I => \N__48020\
        );

    \I__11322\ : ClkMux
    port map (
            O => \N__48396\,
            I => \N__48020\
        );

    \I__11321\ : ClkMux
    port map (
            O => \N__48395\,
            I => \N__48020\
        );

    \I__11320\ : ClkMux
    port map (
            O => \N__48394\,
            I => \N__48020\
        );

    \I__11319\ : ClkMux
    port map (
            O => \N__48393\,
            I => \N__48020\
        );

    \I__11318\ : ClkMux
    port map (
            O => \N__48392\,
            I => \N__48020\
        );

    \I__11317\ : ClkMux
    port map (
            O => \N__48391\,
            I => \N__48020\
        );

    \I__11316\ : ClkMux
    port map (
            O => \N__48390\,
            I => \N__48020\
        );

    \I__11315\ : ClkMux
    port map (
            O => \N__48389\,
            I => \N__48020\
        );

    \I__11314\ : ClkMux
    port map (
            O => \N__48388\,
            I => \N__48020\
        );

    \I__11313\ : ClkMux
    port map (
            O => \N__48387\,
            I => \N__48020\
        );

    \I__11312\ : ClkMux
    port map (
            O => \N__48386\,
            I => \N__48020\
        );

    \I__11311\ : ClkMux
    port map (
            O => \N__48385\,
            I => \N__48020\
        );

    \I__11310\ : ClkMux
    port map (
            O => \N__48384\,
            I => \N__48020\
        );

    \I__11309\ : ClkMux
    port map (
            O => \N__48383\,
            I => \N__48020\
        );

    \I__11308\ : ClkMux
    port map (
            O => \N__48382\,
            I => \N__48020\
        );

    \I__11307\ : ClkMux
    port map (
            O => \N__48381\,
            I => \N__48020\
        );

    \I__11306\ : ClkMux
    port map (
            O => \N__48380\,
            I => \N__48020\
        );

    \I__11305\ : ClkMux
    port map (
            O => \N__48379\,
            I => \N__48020\
        );

    \I__11304\ : ClkMux
    port map (
            O => \N__48378\,
            I => \N__48020\
        );

    \I__11303\ : ClkMux
    port map (
            O => \N__48377\,
            I => \N__48020\
        );

    \I__11302\ : ClkMux
    port map (
            O => \N__48376\,
            I => \N__48020\
        );

    \I__11301\ : ClkMux
    port map (
            O => \N__48375\,
            I => \N__48020\
        );

    \I__11300\ : ClkMux
    port map (
            O => \N__48374\,
            I => \N__48020\
        );

    \I__11299\ : ClkMux
    port map (
            O => \N__48373\,
            I => \N__48020\
        );

    \I__11298\ : ClkMux
    port map (
            O => \N__48372\,
            I => \N__48020\
        );

    \I__11297\ : ClkMux
    port map (
            O => \N__48371\,
            I => \N__48020\
        );

    \I__11296\ : ClkMux
    port map (
            O => \N__48370\,
            I => \N__48020\
        );

    \I__11295\ : ClkMux
    port map (
            O => \N__48369\,
            I => \N__48020\
        );

    \I__11294\ : ClkMux
    port map (
            O => \N__48368\,
            I => \N__48020\
        );

    \I__11293\ : ClkMux
    port map (
            O => \N__48367\,
            I => \N__48020\
        );

    \I__11292\ : ClkMux
    port map (
            O => \N__48366\,
            I => \N__48020\
        );

    \I__11291\ : ClkMux
    port map (
            O => \N__48365\,
            I => \N__48020\
        );

    \I__11290\ : ClkMux
    port map (
            O => \N__48364\,
            I => \N__48020\
        );

    \I__11289\ : ClkMux
    port map (
            O => \N__48363\,
            I => \N__48020\
        );

    \I__11288\ : ClkMux
    port map (
            O => \N__48362\,
            I => \N__48020\
        );

    \I__11287\ : ClkMux
    port map (
            O => \N__48361\,
            I => \N__48020\
        );

    \I__11286\ : ClkMux
    port map (
            O => \N__48360\,
            I => \N__48020\
        );

    \I__11285\ : ClkMux
    port map (
            O => \N__48359\,
            I => \N__48020\
        );

    \I__11284\ : ClkMux
    port map (
            O => \N__48358\,
            I => \N__48020\
        );

    \I__11283\ : ClkMux
    port map (
            O => \N__48357\,
            I => \N__48020\
        );

    \I__11282\ : ClkMux
    port map (
            O => \N__48356\,
            I => \N__48020\
        );

    \I__11281\ : ClkMux
    port map (
            O => \N__48355\,
            I => \N__48020\
        );

    \I__11280\ : ClkMux
    port map (
            O => \N__48354\,
            I => \N__48020\
        );

    \I__11279\ : ClkMux
    port map (
            O => \N__48353\,
            I => \N__48020\
        );

    \I__11278\ : ClkMux
    port map (
            O => \N__48352\,
            I => \N__48020\
        );

    \I__11277\ : ClkMux
    port map (
            O => \N__48351\,
            I => \N__48020\
        );

    \I__11276\ : ClkMux
    port map (
            O => \N__48350\,
            I => \N__48020\
        );

    \I__11275\ : ClkMux
    port map (
            O => \N__48349\,
            I => \N__48020\
        );

    \I__11274\ : ClkMux
    port map (
            O => \N__48348\,
            I => \N__48020\
        );

    \I__11273\ : ClkMux
    port map (
            O => \N__48347\,
            I => \N__48020\
        );

    \I__11272\ : ClkMux
    port map (
            O => \N__48346\,
            I => \N__48020\
        );

    \I__11271\ : ClkMux
    port map (
            O => \N__48345\,
            I => \N__48020\
        );

    \I__11270\ : ClkMux
    port map (
            O => \N__48344\,
            I => \N__48020\
        );

    \I__11269\ : ClkMux
    port map (
            O => \N__48343\,
            I => \N__48020\
        );

    \I__11268\ : ClkMux
    port map (
            O => \N__48342\,
            I => \N__48020\
        );

    \I__11267\ : ClkMux
    port map (
            O => \N__48341\,
            I => \N__48020\
        );

    \I__11266\ : ClkMux
    port map (
            O => \N__48340\,
            I => \N__48020\
        );

    \I__11265\ : ClkMux
    port map (
            O => \N__48339\,
            I => \N__48020\
        );

    \I__11264\ : ClkMux
    port map (
            O => \N__48338\,
            I => \N__48020\
        );

    \I__11263\ : ClkMux
    port map (
            O => \N__48337\,
            I => \N__48020\
        );

    \I__11262\ : ClkMux
    port map (
            O => \N__48336\,
            I => \N__48020\
        );

    \I__11261\ : ClkMux
    port map (
            O => \N__48335\,
            I => \N__48020\
        );

    \I__11260\ : ClkMux
    port map (
            O => \N__48334\,
            I => \N__48020\
        );

    \I__11259\ : ClkMux
    port map (
            O => \N__48333\,
            I => \N__48020\
        );

    \I__11258\ : ClkMux
    port map (
            O => \N__48332\,
            I => \N__48020\
        );

    \I__11257\ : ClkMux
    port map (
            O => \N__48331\,
            I => \N__48020\
        );

    \I__11256\ : ClkMux
    port map (
            O => \N__48330\,
            I => \N__48020\
        );

    \I__11255\ : ClkMux
    port map (
            O => \N__48329\,
            I => \N__48020\
        );

    \I__11254\ : GlobalMux
    port map (
            O => \N__48020\,
            I => clk_100mhz_0
        );

    \I__11253\ : CEMux
    port map (
            O => \N__48017\,
            I => \N__48013\
        );

    \I__11252\ : CEMux
    port map (
            O => \N__48016\,
            I => \N__48009\
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__48013\,
            I => \N__48005\
        );

    \I__11250\ : CEMux
    port map (
            O => \N__48012\,
            I => \N__48002\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__48009\,
            I => \N__47999\
        );

    \I__11248\ : CEMux
    port map (
            O => \N__48008\,
            I => \N__47996\
        );

    \I__11247\ : Span4Mux_v
    port map (
            O => \N__48005\,
            I => \N__47989\
        );

    \I__11246\ : LocalMux
    port map (
            O => \N__48002\,
            I => \N__47989\
        );

    \I__11245\ : Span4Mux_h
    port map (
            O => \N__47999\,
            I => \N__47982\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__47996\,
            I => \N__47982\
        );

    \I__11243\ : CEMux
    port map (
            O => \N__47995\,
            I => \N__47979\
        );

    \I__11242\ : CEMux
    port map (
            O => \N__47994\,
            I => \N__47976\
        );

    \I__11241\ : Span4Mux_v
    port map (
            O => \N__47989\,
            I => \N__47973\
        );

    \I__11240\ : CEMux
    port map (
            O => \N__47988\,
            I => \N__47970\
        );

    \I__11239\ : CEMux
    port map (
            O => \N__47987\,
            I => \N__47967\
        );

    \I__11238\ : Span4Mux_h
    port map (
            O => \N__47982\,
            I => \N__47960\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__47979\,
            I => \N__47960\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__47976\,
            I => \N__47960\
        );

    \I__11235\ : Span4Mux_h
    port map (
            O => \N__47973\,
            I => \N__47955\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__47970\,
            I => \N__47955\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__47967\,
            I => \N__47951\
        );

    \I__11232\ : Span4Mux_v
    port map (
            O => \N__47960\,
            I => \N__47948\
        );

    \I__11231\ : Span4Mux_h
    port map (
            O => \N__47955\,
            I => \N__47945\
        );

    \I__11230\ : CEMux
    port map (
            O => \N__47954\,
            I => \N__47942\
        );

    \I__11229\ : Span4Mux_v
    port map (
            O => \N__47951\,
            I => \N__47937\
        );

    \I__11228\ : Span4Mux_h
    port map (
            O => \N__47948\,
            I => \N__47937\
        );

    \I__11227\ : Span4Mux_v
    port map (
            O => \N__47945\,
            I => \N__47932\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__47942\,
            I => \N__47932\
        );

    \I__11225\ : Odrv4
    port map (
            O => \N__47937\,
            I => \current_shift_inst.timer_s1.N_180_i_g\
        );

    \I__11224\ : Odrv4
    port map (
            O => \N__47932\,
            I => \current_shift_inst.timer_s1.N_180_i_g\
        );

    \I__11223\ : CascadeMux
    port map (
            O => \N__47927\,
            I => \N__47919\
        );

    \I__11222\ : CascadeMux
    port map (
            O => \N__47926\,
            I => \N__47915\
        );

    \I__11221\ : InMux
    port map (
            O => \N__47925\,
            I => \N__47912\
        );

    \I__11220\ : InMux
    port map (
            O => \N__47924\,
            I => \N__47909\
        );

    \I__11219\ : InMux
    port map (
            O => \N__47923\,
            I => \N__47906\
        );

    \I__11218\ : InMux
    port map (
            O => \N__47922\,
            I => \N__47903\
        );

    \I__11217\ : InMux
    port map (
            O => \N__47919\,
            I => \N__47900\
        );

    \I__11216\ : InMux
    port map (
            O => \N__47918\,
            I => \N__47897\
        );

    \I__11215\ : InMux
    port map (
            O => \N__47915\,
            I => \N__47894\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__47912\,
            I => \N__47891\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__47909\,
            I => \N__47888\
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__47906\,
            I => \N__47885\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__47903\,
            I => \N__47844\
        );

    \I__11210\ : LocalMux
    port map (
            O => \N__47900\,
            I => \N__47781\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__47897\,
            I => \N__47762\
        );

    \I__11208\ : LocalMux
    port map (
            O => \N__47894\,
            I => \N__47743\
        );

    \I__11207\ : Glb2LocalMux
    port map (
            O => \N__47891\,
            I => \N__47444\
        );

    \I__11206\ : Glb2LocalMux
    port map (
            O => \N__47888\,
            I => \N__47444\
        );

    \I__11205\ : Glb2LocalMux
    port map (
            O => \N__47885\,
            I => \N__47444\
        );

    \I__11204\ : SRMux
    port map (
            O => \N__47884\,
            I => \N__47444\
        );

    \I__11203\ : SRMux
    port map (
            O => \N__47883\,
            I => \N__47444\
        );

    \I__11202\ : SRMux
    port map (
            O => \N__47882\,
            I => \N__47444\
        );

    \I__11201\ : SRMux
    port map (
            O => \N__47881\,
            I => \N__47444\
        );

    \I__11200\ : SRMux
    port map (
            O => \N__47880\,
            I => \N__47444\
        );

    \I__11199\ : SRMux
    port map (
            O => \N__47879\,
            I => \N__47444\
        );

    \I__11198\ : SRMux
    port map (
            O => \N__47878\,
            I => \N__47444\
        );

    \I__11197\ : SRMux
    port map (
            O => \N__47877\,
            I => \N__47444\
        );

    \I__11196\ : SRMux
    port map (
            O => \N__47876\,
            I => \N__47444\
        );

    \I__11195\ : SRMux
    port map (
            O => \N__47875\,
            I => \N__47444\
        );

    \I__11194\ : SRMux
    port map (
            O => \N__47874\,
            I => \N__47444\
        );

    \I__11193\ : SRMux
    port map (
            O => \N__47873\,
            I => \N__47444\
        );

    \I__11192\ : SRMux
    port map (
            O => \N__47872\,
            I => \N__47444\
        );

    \I__11191\ : SRMux
    port map (
            O => \N__47871\,
            I => \N__47444\
        );

    \I__11190\ : SRMux
    port map (
            O => \N__47870\,
            I => \N__47444\
        );

    \I__11189\ : SRMux
    port map (
            O => \N__47869\,
            I => \N__47444\
        );

    \I__11188\ : SRMux
    port map (
            O => \N__47868\,
            I => \N__47444\
        );

    \I__11187\ : SRMux
    port map (
            O => \N__47867\,
            I => \N__47444\
        );

    \I__11186\ : SRMux
    port map (
            O => \N__47866\,
            I => \N__47444\
        );

    \I__11185\ : SRMux
    port map (
            O => \N__47865\,
            I => \N__47444\
        );

    \I__11184\ : SRMux
    port map (
            O => \N__47864\,
            I => \N__47444\
        );

    \I__11183\ : SRMux
    port map (
            O => \N__47863\,
            I => \N__47444\
        );

    \I__11182\ : SRMux
    port map (
            O => \N__47862\,
            I => \N__47444\
        );

    \I__11181\ : SRMux
    port map (
            O => \N__47861\,
            I => \N__47444\
        );

    \I__11180\ : SRMux
    port map (
            O => \N__47860\,
            I => \N__47444\
        );

    \I__11179\ : SRMux
    port map (
            O => \N__47859\,
            I => \N__47444\
        );

    \I__11178\ : SRMux
    port map (
            O => \N__47858\,
            I => \N__47444\
        );

    \I__11177\ : SRMux
    port map (
            O => \N__47857\,
            I => \N__47444\
        );

    \I__11176\ : SRMux
    port map (
            O => \N__47856\,
            I => \N__47444\
        );

    \I__11175\ : SRMux
    port map (
            O => \N__47855\,
            I => \N__47444\
        );

    \I__11174\ : SRMux
    port map (
            O => \N__47854\,
            I => \N__47444\
        );

    \I__11173\ : SRMux
    port map (
            O => \N__47853\,
            I => \N__47444\
        );

    \I__11172\ : SRMux
    port map (
            O => \N__47852\,
            I => \N__47444\
        );

    \I__11171\ : SRMux
    port map (
            O => \N__47851\,
            I => \N__47444\
        );

    \I__11170\ : SRMux
    port map (
            O => \N__47850\,
            I => \N__47444\
        );

    \I__11169\ : SRMux
    port map (
            O => \N__47849\,
            I => \N__47444\
        );

    \I__11168\ : SRMux
    port map (
            O => \N__47848\,
            I => \N__47444\
        );

    \I__11167\ : SRMux
    port map (
            O => \N__47847\,
            I => \N__47444\
        );

    \I__11166\ : Glb2LocalMux
    port map (
            O => \N__47844\,
            I => \N__47444\
        );

    \I__11165\ : SRMux
    port map (
            O => \N__47843\,
            I => \N__47444\
        );

    \I__11164\ : SRMux
    port map (
            O => \N__47842\,
            I => \N__47444\
        );

    \I__11163\ : SRMux
    port map (
            O => \N__47841\,
            I => \N__47444\
        );

    \I__11162\ : SRMux
    port map (
            O => \N__47840\,
            I => \N__47444\
        );

    \I__11161\ : SRMux
    port map (
            O => \N__47839\,
            I => \N__47444\
        );

    \I__11160\ : SRMux
    port map (
            O => \N__47838\,
            I => \N__47444\
        );

    \I__11159\ : SRMux
    port map (
            O => \N__47837\,
            I => \N__47444\
        );

    \I__11158\ : SRMux
    port map (
            O => \N__47836\,
            I => \N__47444\
        );

    \I__11157\ : SRMux
    port map (
            O => \N__47835\,
            I => \N__47444\
        );

    \I__11156\ : SRMux
    port map (
            O => \N__47834\,
            I => \N__47444\
        );

    \I__11155\ : SRMux
    port map (
            O => \N__47833\,
            I => \N__47444\
        );

    \I__11154\ : SRMux
    port map (
            O => \N__47832\,
            I => \N__47444\
        );

    \I__11153\ : SRMux
    port map (
            O => \N__47831\,
            I => \N__47444\
        );

    \I__11152\ : SRMux
    port map (
            O => \N__47830\,
            I => \N__47444\
        );

    \I__11151\ : SRMux
    port map (
            O => \N__47829\,
            I => \N__47444\
        );

    \I__11150\ : SRMux
    port map (
            O => \N__47828\,
            I => \N__47444\
        );

    \I__11149\ : SRMux
    port map (
            O => \N__47827\,
            I => \N__47444\
        );

    \I__11148\ : SRMux
    port map (
            O => \N__47826\,
            I => \N__47444\
        );

    \I__11147\ : SRMux
    port map (
            O => \N__47825\,
            I => \N__47444\
        );

    \I__11146\ : SRMux
    port map (
            O => \N__47824\,
            I => \N__47444\
        );

    \I__11145\ : SRMux
    port map (
            O => \N__47823\,
            I => \N__47444\
        );

    \I__11144\ : SRMux
    port map (
            O => \N__47822\,
            I => \N__47444\
        );

    \I__11143\ : SRMux
    port map (
            O => \N__47821\,
            I => \N__47444\
        );

    \I__11142\ : SRMux
    port map (
            O => \N__47820\,
            I => \N__47444\
        );

    \I__11141\ : SRMux
    port map (
            O => \N__47819\,
            I => \N__47444\
        );

    \I__11140\ : SRMux
    port map (
            O => \N__47818\,
            I => \N__47444\
        );

    \I__11139\ : SRMux
    port map (
            O => \N__47817\,
            I => \N__47444\
        );

    \I__11138\ : SRMux
    port map (
            O => \N__47816\,
            I => \N__47444\
        );

    \I__11137\ : SRMux
    port map (
            O => \N__47815\,
            I => \N__47444\
        );

    \I__11136\ : SRMux
    port map (
            O => \N__47814\,
            I => \N__47444\
        );

    \I__11135\ : SRMux
    port map (
            O => \N__47813\,
            I => \N__47444\
        );

    \I__11134\ : SRMux
    port map (
            O => \N__47812\,
            I => \N__47444\
        );

    \I__11133\ : SRMux
    port map (
            O => \N__47811\,
            I => \N__47444\
        );

    \I__11132\ : SRMux
    port map (
            O => \N__47810\,
            I => \N__47444\
        );

    \I__11131\ : SRMux
    port map (
            O => \N__47809\,
            I => \N__47444\
        );

    \I__11130\ : SRMux
    port map (
            O => \N__47808\,
            I => \N__47444\
        );

    \I__11129\ : SRMux
    port map (
            O => \N__47807\,
            I => \N__47444\
        );

    \I__11128\ : SRMux
    port map (
            O => \N__47806\,
            I => \N__47444\
        );

    \I__11127\ : SRMux
    port map (
            O => \N__47805\,
            I => \N__47444\
        );

    \I__11126\ : SRMux
    port map (
            O => \N__47804\,
            I => \N__47444\
        );

    \I__11125\ : SRMux
    port map (
            O => \N__47803\,
            I => \N__47444\
        );

    \I__11124\ : SRMux
    port map (
            O => \N__47802\,
            I => \N__47444\
        );

    \I__11123\ : SRMux
    port map (
            O => \N__47801\,
            I => \N__47444\
        );

    \I__11122\ : SRMux
    port map (
            O => \N__47800\,
            I => \N__47444\
        );

    \I__11121\ : SRMux
    port map (
            O => \N__47799\,
            I => \N__47444\
        );

    \I__11120\ : SRMux
    port map (
            O => \N__47798\,
            I => \N__47444\
        );

    \I__11119\ : SRMux
    port map (
            O => \N__47797\,
            I => \N__47444\
        );

    \I__11118\ : SRMux
    port map (
            O => \N__47796\,
            I => \N__47444\
        );

    \I__11117\ : SRMux
    port map (
            O => \N__47795\,
            I => \N__47444\
        );

    \I__11116\ : SRMux
    port map (
            O => \N__47794\,
            I => \N__47444\
        );

    \I__11115\ : SRMux
    port map (
            O => \N__47793\,
            I => \N__47444\
        );

    \I__11114\ : SRMux
    port map (
            O => \N__47792\,
            I => \N__47444\
        );

    \I__11113\ : SRMux
    port map (
            O => \N__47791\,
            I => \N__47444\
        );

    \I__11112\ : SRMux
    port map (
            O => \N__47790\,
            I => \N__47444\
        );

    \I__11111\ : SRMux
    port map (
            O => \N__47789\,
            I => \N__47444\
        );

    \I__11110\ : SRMux
    port map (
            O => \N__47788\,
            I => \N__47444\
        );

    \I__11109\ : SRMux
    port map (
            O => \N__47787\,
            I => \N__47444\
        );

    \I__11108\ : SRMux
    port map (
            O => \N__47786\,
            I => \N__47444\
        );

    \I__11107\ : SRMux
    port map (
            O => \N__47785\,
            I => \N__47444\
        );

    \I__11106\ : SRMux
    port map (
            O => \N__47784\,
            I => \N__47444\
        );

    \I__11105\ : Glb2LocalMux
    port map (
            O => \N__47781\,
            I => \N__47444\
        );

    \I__11104\ : SRMux
    port map (
            O => \N__47780\,
            I => \N__47444\
        );

    \I__11103\ : SRMux
    port map (
            O => \N__47779\,
            I => \N__47444\
        );

    \I__11102\ : SRMux
    port map (
            O => \N__47778\,
            I => \N__47444\
        );

    \I__11101\ : SRMux
    port map (
            O => \N__47777\,
            I => \N__47444\
        );

    \I__11100\ : SRMux
    port map (
            O => \N__47776\,
            I => \N__47444\
        );

    \I__11099\ : SRMux
    port map (
            O => \N__47775\,
            I => \N__47444\
        );

    \I__11098\ : SRMux
    port map (
            O => \N__47774\,
            I => \N__47444\
        );

    \I__11097\ : SRMux
    port map (
            O => \N__47773\,
            I => \N__47444\
        );

    \I__11096\ : SRMux
    port map (
            O => \N__47772\,
            I => \N__47444\
        );

    \I__11095\ : SRMux
    port map (
            O => \N__47771\,
            I => \N__47444\
        );

    \I__11094\ : SRMux
    port map (
            O => \N__47770\,
            I => \N__47444\
        );

    \I__11093\ : SRMux
    port map (
            O => \N__47769\,
            I => \N__47444\
        );

    \I__11092\ : SRMux
    port map (
            O => \N__47768\,
            I => \N__47444\
        );

    \I__11091\ : SRMux
    port map (
            O => \N__47767\,
            I => \N__47444\
        );

    \I__11090\ : SRMux
    port map (
            O => \N__47766\,
            I => \N__47444\
        );

    \I__11089\ : SRMux
    port map (
            O => \N__47765\,
            I => \N__47444\
        );

    \I__11088\ : Glb2LocalMux
    port map (
            O => \N__47762\,
            I => \N__47444\
        );

    \I__11087\ : SRMux
    port map (
            O => \N__47761\,
            I => \N__47444\
        );

    \I__11086\ : SRMux
    port map (
            O => \N__47760\,
            I => \N__47444\
        );

    \I__11085\ : SRMux
    port map (
            O => \N__47759\,
            I => \N__47444\
        );

    \I__11084\ : SRMux
    port map (
            O => \N__47758\,
            I => \N__47444\
        );

    \I__11083\ : SRMux
    port map (
            O => \N__47757\,
            I => \N__47444\
        );

    \I__11082\ : SRMux
    port map (
            O => \N__47756\,
            I => \N__47444\
        );

    \I__11081\ : SRMux
    port map (
            O => \N__47755\,
            I => \N__47444\
        );

    \I__11080\ : SRMux
    port map (
            O => \N__47754\,
            I => \N__47444\
        );

    \I__11079\ : SRMux
    port map (
            O => \N__47753\,
            I => \N__47444\
        );

    \I__11078\ : SRMux
    port map (
            O => \N__47752\,
            I => \N__47444\
        );

    \I__11077\ : SRMux
    port map (
            O => \N__47751\,
            I => \N__47444\
        );

    \I__11076\ : SRMux
    port map (
            O => \N__47750\,
            I => \N__47444\
        );

    \I__11075\ : SRMux
    port map (
            O => \N__47749\,
            I => \N__47444\
        );

    \I__11074\ : SRMux
    port map (
            O => \N__47748\,
            I => \N__47444\
        );

    \I__11073\ : SRMux
    port map (
            O => \N__47747\,
            I => \N__47444\
        );

    \I__11072\ : SRMux
    port map (
            O => \N__47746\,
            I => \N__47444\
        );

    \I__11071\ : Glb2LocalMux
    port map (
            O => \N__47743\,
            I => \N__47444\
        );

    \I__11070\ : SRMux
    port map (
            O => \N__47742\,
            I => \N__47444\
        );

    \I__11069\ : SRMux
    port map (
            O => \N__47741\,
            I => \N__47444\
        );

    \I__11068\ : SRMux
    port map (
            O => \N__47740\,
            I => \N__47444\
        );

    \I__11067\ : SRMux
    port map (
            O => \N__47739\,
            I => \N__47444\
        );

    \I__11066\ : SRMux
    port map (
            O => \N__47738\,
            I => \N__47444\
        );

    \I__11065\ : SRMux
    port map (
            O => \N__47737\,
            I => \N__47444\
        );

    \I__11064\ : SRMux
    port map (
            O => \N__47736\,
            I => \N__47444\
        );

    \I__11063\ : SRMux
    port map (
            O => \N__47735\,
            I => \N__47444\
        );

    \I__11062\ : GlobalMux
    port map (
            O => \N__47444\,
            I => \N__47441\
        );

    \I__11061\ : gio2CtrlBuf
    port map (
            O => \N__47441\,
            I => red_c_g
        );

    \I__11060\ : CascadeMux
    port map (
            O => \N__47438\,
            I => \N__47434\
        );

    \I__11059\ : InMux
    port map (
            O => \N__47437\,
            I => \N__47431\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47434\,
            I => \N__47428\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__47431\,
            I => \N__47423\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__47428\,
            I => \N__47420\
        );

    \I__11055\ : InMux
    port map (
            O => \N__47427\,
            I => \N__47417\
        );

    \I__11054\ : InMux
    port map (
            O => \N__47426\,
            I => \N__47414\
        );

    \I__11053\ : Span4Mux_h
    port map (
            O => \N__47423\,
            I => \N__47411\
        );

    \I__11052\ : Span4Mux_v
    port map (
            O => \N__47420\,
            I => \N__47408\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__47417\,
            I => \N__47403\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__47414\,
            I => \N__47403\
        );

    \I__11049\ : Span4Mux_v
    port map (
            O => \N__47411\,
            I => \N__47398\
        );

    \I__11048\ : Span4Mux_v
    port map (
            O => \N__47408\,
            I => \N__47398\
        );

    \I__11047\ : Span4Mux_h
    port map (
            O => \N__47403\,
            I => \N__47395\
        );

    \I__11046\ : Odrv4
    port map (
            O => \N__47398\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__11045\ : Odrv4
    port map (
            O => \N__47395\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__11044\ : InMux
    port map (
            O => \N__47390\,
            I => \N__47387\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__47387\,
            I => \N__47382\
        );

    \I__11042\ : InMux
    port map (
            O => \N__47386\,
            I => \N__47379\
        );

    \I__11041\ : InMux
    port map (
            O => \N__47385\,
            I => \N__47376\
        );

    \I__11040\ : Odrv4
    port map (
            O => \N__47382\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__47379\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__47376\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__11037\ : InMux
    port map (
            O => \N__47369\,
            I => \N__47366\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__47366\,
            I => \N__47363\
        );

    \I__11035\ : Span4Mux_v
    port map (
            O => \N__47363\,
            I => \N__47360\
        );

    \I__11034\ : Odrv4
    port map (
            O => \N__47360\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__11033\ : InMux
    port map (
            O => \N__47357\,
            I => \N__47353\
        );

    \I__11032\ : InMux
    port map (
            O => \N__47356\,
            I => \N__47350\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__47353\,
            I => \N__47346\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__47350\,
            I => \N__47343\
        );

    \I__11029\ : InMux
    port map (
            O => \N__47349\,
            I => \N__47340\
        );

    \I__11028\ : Span4Mux_v
    port map (
            O => \N__47346\,
            I => \N__47337\
        );

    \I__11027\ : Span4Mux_v
    port map (
            O => \N__47343\,
            I => \N__47331\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__47340\,
            I => \N__47331\
        );

    \I__11025\ : Span4Mux_h
    port map (
            O => \N__47337\,
            I => \N__47328\
        );

    \I__11024\ : InMux
    port map (
            O => \N__47336\,
            I => \N__47325\
        );

    \I__11023\ : Odrv4
    port map (
            O => \N__47331\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11022\ : Odrv4
    port map (
            O => \N__47328\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__47325\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__11020\ : CascadeMux
    port map (
            O => \N__47318\,
            I => \N__47314\
        );

    \I__11019\ : InMux
    port map (
            O => \N__47317\,
            I => \N__47310\
        );

    \I__11018\ : InMux
    port map (
            O => \N__47314\,
            I => \N__47307\
        );

    \I__11017\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47304\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__47310\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__47307\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__11014\ : LocalMux
    port map (
            O => \N__47304\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__11013\ : InMux
    port map (
            O => \N__47297\,
            I => \N__47294\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__47294\,
            I => \N__47291\
        );

    \I__11011\ : Odrv4
    port map (
            O => \N__47291\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__11010\ : InMux
    port map (
            O => \N__47288\,
            I => \N__47283\
        );

    \I__11009\ : InMux
    port map (
            O => \N__47287\,
            I => \N__47277\
        );

    \I__11008\ : InMux
    port map (
            O => \N__47286\,
            I => \N__47277\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__47283\,
            I => \N__47274\
        );

    \I__11006\ : InMux
    port map (
            O => \N__47282\,
            I => \N__47271\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__47277\,
            I => \N__47268\
        );

    \I__11004\ : Span4Mux_h
    port map (
            O => \N__47274\,
            I => \N__47265\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__47271\,
            I => \N__47260\
        );

    \I__11002\ : Span4Mux_h
    port map (
            O => \N__47268\,
            I => \N__47260\
        );

    \I__11001\ : Odrv4
    port map (
            O => \N__47265\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__11000\ : Odrv4
    port map (
            O => \N__47260\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__10999\ : InMux
    port map (
            O => \N__47255\,
            I => \N__47250\
        );

    \I__10998\ : InMux
    port map (
            O => \N__47254\,
            I => \N__47247\
        );

    \I__10997\ : InMux
    port map (
            O => \N__47253\,
            I => \N__47244\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__47250\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__47247\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10994\ : LocalMux
    port map (
            O => \N__47244\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__10993\ : InMux
    port map (
            O => \N__47237\,
            I => \N__47234\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__47234\,
            I => \N__47231\
        );

    \I__10991\ : Odrv12
    port map (
            O => \N__47231\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__10990\ : CascadeMux
    port map (
            O => \N__47228\,
            I => \N__47224\
        );

    \I__10989\ : InMux
    port map (
            O => \N__47227\,
            I => \N__47220\
        );

    \I__10988\ : InMux
    port map (
            O => \N__47224\,
            I => \N__47217\
        );

    \I__10987\ : InMux
    port map (
            O => \N__47223\,
            I => \N__47214\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__47220\,
            I => \N__47211\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__47217\,
            I => \N__47206\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__47214\,
            I => \N__47206\
        );

    \I__10983\ : Span4Mux_h
    port map (
            O => \N__47211\,
            I => \N__47202\
        );

    \I__10982\ : Span4Mux_v
    port map (
            O => \N__47206\,
            I => \N__47199\
        );

    \I__10981\ : InMux
    port map (
            O => \N__47205\,
            I => \N__47196\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__47202\,
            I => \N__47189\
        );

    \I__10979\ : Span4Mux_v
    port map (
            O => \N__47199\,
            I => \N__47189\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__47196\,
            I => \N__47189\
        );

    \I__10977\ : Odrv4
    port map (
            O => \N__47189\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__10976\ : InMux
    port map (
            O => \N__47186\,
            I => \N__47181\
        );

    \I__10975\ : InMux
    port map (
            O => \N__47185\,
            I => \N__47178\
        );

    \I__10974\ : InMux
    port map (
            O => \N__47184\,
            I => \N__47175\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__47181\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__47178\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__47175\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__10970\ : InMux
    port map (
            O => \N__47168\,
            I => \N__47165\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__47165\,
            I => \N__47162\
        );

    \I__10968\ : Odrv4
    port map (
            O => \N__47162\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__10967\ : InMux
    port map (
            O => \N__47159\,
            I => \N__47155\
        );

    \I__10966\ : InMux
    port map (
            O => \N__47158\,
            I => \N__47152\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__47155\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__47152\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__10963\ : InMux
    port map (
            O => \N__47147\,
            I => \N__47144\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__47144\,
            I => \N__47141\
        );

    \I__10961\ : Odrv4
    port map (
            O => \N__47141\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__10960\ : InMux
    port map (
            O => \N__47138\,
            I => \N__47133\
        );

    \I__10959\ : InMux
    port map (
            O => \N__47137\,
            I => \N__47130\
        );

    \I__10958\ : InMux
    port map (
            O => \N__47136\,
            I => \N__47127\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__47133\,
            I => \N__47124\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__47130\,
            I => \N__47121\
        );

    \I__10955\ : LocalMux
    port map (
            O => \N__47127\,
            I => \N__47116\
        );

    \I__10954\ : Span4Mux_v
    port map (
            O => \N__47124\,
            I => \N__47116\
        );

    \I__10953\ : Span4Mux_v
    port map (
            O => \N__47121\,
            I => \N__47110\
        );

    \I__10952\ : Span4Mux_h
    port map (
            O => \N__47116\,
            I => \N__47110\
        );

    \I__10951\ : InMux
    port map (
            O => \N__47115\,
            I => \N__47107\
        );

    \I__10950\ : Odrv4
    port map (
            O => \N__47110\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__47107\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__10948\ : InMux
    port map (
            O => \N__47102\,
            I => \N__47099\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__47099\,
            I => \N__47096\
        );

    \I__10946\ : Span4Mux_v
    port map (
            O => \N__47096\,
            I => \N__47091\
        );

    \I__10945\ : InMux
    port map (
            O => \N__47095\,
            I => \N__47088\
        );

    \I__10944\ : InMux
    port map (
            O => \N__47094\,
            I => \N__47085\
        );

    \I__10943\ : Odrv4
    port map (
            O => \N__47091\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__47088\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__47085\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__10940\ : InMux
    port map (
            O => \N__47078\,
            I => \N__47075\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__47075\,
            I => \N__47072\
        );

    \I__10938\ : Odrv12
    port map (
            O => \N__47072\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__10937\ : InMux
    port map (
            O => \N__47069\,
            I => \N__47063\
        );

    \I__10936\ : InMux
    port map (
            O => \N__47068\,
            I => \N__47060\
        );

    \I__10935\ : InMux
    port map (
            O => \N__47067\,
            I => \N__47057\
        );

    \I__10934\ : InMux
    port map (
            O => \N__47066\,
            I => \N__47054\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__47063\,
            I => \N__47051\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__47060\,
            I => \N__47048\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__47057\,
            I => \N__47045\
        );

    \I__10930\ : LocalMux
    port map (
            O => \N__47054\,
            I => \N__47042\
        );

    \I__10929\ : Span12Mux_v
    port map (
            O => \N__47051\,
            I => \N__47037\
        );

    \I__10928\ : Span12Mux_s10_h
    port map (
            O => \N__47048\,
            I => \N__47037\
        );

    \I__10927\ : Span4Mux_v
    port map (
            O => \N__47045\,
            I => \N__47034\
        );

    \I__10926\ : Odrv4
    port map (
            O => \N__47042\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__10925\ : Odrv12
    port map (
            O => \N__47037\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__10924\ : Odrv4
    port map (
            O => \N__47034\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__10923\ : InMux
    port map (
            O => \N__47027\,
            I => \N__47024\
        );

    \I__10922\ : LocalMux
    port map (
            O => \N__47024\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47021\,
            I => \N__47018\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__47018\,
            I => \N__47015\
        );

    \I__10919\ : Span4Mux_h
    port map (
            O => \N__47015\,
            I => \N__47012\
        );

    \I__10918\ : Odrv4
    port map (
            O => \N__47012\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__10917\ : CascadeMux
    port map (
            O => \N__47009\,
            I => \N__47005\
        );

    \I__10916\ : InMux
    port map (
            O => \N__47008\,
            I => \N__47001\
        );

    \I__10915\ : InMux
    port map (
            O => \N__47005\,
            I => \N__46996\
        );

    \I__10914\ : InMux
    port map (
            O => \N__47004\,
            I => \N__46996\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__47001\,
            I => \N__46991\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__46996\,
            I => \N__46991\
        );

    \I__10911\ : Span4Mux_h
    port map (
            O => \N__46991\,
            I => \N__46987\
        );

    \I__10910\ : InMux
    port map (
            O => \N__46990\,
            I => \N__46984\
        );

    \I__10909\ : Odrv4
    port map (
            O => \N__46987\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__46984\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__10907\ : InMux
    port map (
            O => \N__46979\,
            I => \N__46974\
        );

    \I__10906\ : InMux
    port map (
            O => \N__46978\,
            I => \N__46969\
        );

    \I__10905\ : InMux
    port map (
            O => \N__46977\,
            I => \N__46969\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__46974\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__46969\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__10902\ : InMux
    port map (
            O => \N__46964\,
            I => \N__46956\
        );

    \I__10901\ : InMux
    port map (
            O => \N__46963\,
            I => \N__46956\
        );

    \I__10900\ : InMux
    port map (
            O => \N__46962\,
            I => \N__46951\
        );

    \I__10899\ : InMux
    port map (
            O => \N__46961\,
            I => \N__46951\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__46956\,
            I => \N__46948\
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__46951\,
            I => \N__46945\
        );

    \I__10896\ : Span4Mux_h
    port map (
            O => \N__46948\,
            I => \N__46942\
        );

    \I__10895\ : Odrv4
    port map (
            O => \N__46945\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10894\ : Odrv4
    port map (
            O => \N__46942\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10893\ : InMux
    port map (
            O => \N__46937\,
            I => \N__46934\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__46934\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__10891\ : CascadeMux
    port map (
            O => \N__46931\,
            I => \N__46927\
        );

    \I__10890\ : InMux
    port map (
            O => \N__46930\,
            I => \N__46923\
        );

    \I__10889\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46920\
        );

    \I__10888\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46917\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__46923\,
            I => \N__46914\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__46920\,
            I => \N__46911\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__46917\,
            I => \N__46908\
        );

    \I__10884\ : Span4Mux_v
    port map (
            O => \N__46914\,
            I => \N__46905\
        );

    \I__10883\ : Span4Mux_v
    port map (
            O => \N__46911\,
            I => \N__46901\
        );

    \I__10882\ : Span4Mux_h
    port map (
            O => \N__46908\,
            I => \N__46896\
        );

    \I__10881\ : Span4Mux_h
    port map (
            O => \N__46905\,
            I => \N__46896\
        );

    \I__10880\ : InMux
    port map (
            O => \N__46904\,
            I => \N__46893\
        );

    \I__10879\ : Odrv4
    port map (
            O => \N__46901\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10878\ : Odrv4
    port map (
            O => \N__46896\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__46893\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46886\,
            I => \N__46883\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__46883\,
            I => \N__46878\
        );

    \I__10874\ : InMux
    port map (
            O => \N__46882\,
            I => \N__46875\
        );

    \I__10873\ : InMux
    port map (
            O => \N__46881\,
            I => \N__46872\
        );

    \I__10872\ : Odrv4
    port map (
            O => \N__46878\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__46875\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__46872\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__10869\ : InMux
    port map (
            O => \N__46865\,
            I => \N__46862\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__46862\,
            I => \N__46859\
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__46859\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__10866\ : InMux
    port map (
            O => \N__46856\,
            I => \N__46851\
        );

    \I__10865\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46848\
        );

    \I__10864\ : InMux
    port map (
            O => \N__46854\,
            I => \N__46845\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__46851\,
            I => \N__46842\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__46848\,
            I => \N__46839\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__46845\,
            I => \N__46836\
        );

    \I__10860\ : Span4Mux_v
    port map (
            O => \N__46842\,
            I => \N__46833\
        );

    \I__10859\ : Span4Mux_v
    port map (
            O => \N__46839\,
            I => \N__46829\
        );

    \I__10858\ : Span4Mux_v
    port map (
            O => \N__46836\,
            I => \N__46824\
        );

    \I__10857\ : Span4Mux_h
    port map (
            O => \N__46833\,
            I => \N__46824\
        );

    \I__10856\ : InMux
    port map (
            O => \N__46832\,
            I => \N__46821\
        );

    \I__10855\ : Odrv4
    port map (
            O => \N__46829\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__10854\ : Odrv4
    port map (
            O => \N__46824\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__46821\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__10852\ : InMux
    port map (
            O => \N__46814\,
            I => \N__46811\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__46811\,
            I => \N__46806\
        );

    \I__10850\ : InMux
    port map (
            O => \N__46810\,
            I => \N__46803\
        );

    \I__10849\ : InMux
    port map (
            O => \N__46809\,
            I => \N__46800\
        );

    \I__10848\ : Odrv12
    port map (
            O => \N__46806\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__46803\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__10846\ : LocalMux
    port map (
            O => \N__46800\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46793\,
            I => \N__46790\
        );

    \I__10844\ : LocalMux
    port map (
            O => \N__46790\,
            I => \N__46787\
        );

    \I__10843\ : Odrv4
    port map (
            O => \N__46787\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__10842\ : CascadeMux
    port map (
            O => \N__46784\,
            I => \N__46779\
        );

    \I__10841\ : CascadeMux
    port map (
            O => \N__46783\,
            I => \N__46776\
        );

    \I__10840\ : InMux
    port map (
            O => \N__46782\,
            I => \N__46773\
        );

    \I__10839\ : InMux
    port map (
            O => \N__46779\,
            I => \N__46770\
        );

    \I__10838\ : InMux
    port map (
            O => \N__46776\,
            I => \N__46767\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__46773\,
            I => \N__46764\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__46770\,
            I => \N__46761\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__46767\,
            I => \N__46758\
        );

    \I__10834\ : Span4Mux_h
    port map (
            O => \N__46764\,
            I => \N__46755\
        );

    \I__10833\ : Span4Mux_h
    port map (
            O => \N__46761\,
            I => \N__46751\
        );

    \I__10832\ : Span4Mux_v
    port map (
            O => \N__46758\,
            I => \N__46746\
        );

    \I__10831\ : Span4Mux_v
    port map (
            O => \N__46755\,
            I => \N__46746\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46754\,
            I => \N__46743\
        );

    \I__10829\ : Odrv4
    port map (
            O => \N__46751\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10828\ : Odrv4
    port map (
            O => \N__46746\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__46743\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10826\ : InMux
    port map (
            O => \N__46736\,
            I => \N__46733\
        );

    \I__10825\ : LocalMux
    port map (
            O => \N__46733\,
            I => \N__46728\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46732\,
            I => \N__46725\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46731\,
            I => \N__46722\
        );

    \I__10822\ : Odrv12
    port map (
            O => \N__46728\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__46725\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__46722\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10819\ : InMux
    port map (
            O => \N__46715\,
            I => \N__46712\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__46712\,
            I => \N__46709\
        );

    \I__10817\ : Odrv4
    port map (
            O => \N__46709\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__10816\ : CascadeMux
    port map (
            O => \N__46706\,
            I => \N__46703\
        );

    \I__10815\ : InMux
    port map (
            O => \N__46703\,
            I => \N__46698\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46702\,
            I => \N__46695\
        );

    \I__10813\ : InMux
    port map (
            O => \N__46701\,
            I => \N__46691\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__46698\,
            I => \N__46688\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__46695\,
            I => \N__46685\
        );

    \I__10810\ : InMux
    port map (
            O => \N__46694\,
            I => \N__46682\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__46691\,
            I => \N__46679\
        );

    \I__10808\ : Span4Mux_h
    port map (
            O => \N__46688\,
            I => \N__46676\
        );

    \I__10807\ : Span4Mux_v
    port map (
            O => \N__46685\,
            I => \N__46673\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__46682\,
            I => \N__46670\
        );

    \I__10805\ : Span4Mux_h
    port map (
            O => \N__46679\,
            I => \N__46667\
        );

    \I__10804\ : Span4Mux_v
    port map (
            O => \N__46676\,
            I => \N__46664\
        );

    \I__10803\ : Span4Mux_h
    port map (
            O => \N__46673\,
            I => \N__46661\
        );

    \I__10802\ : Span12Mux_v
    port map (
            O => \N__46670\,
            I => \N__46658\
        );

    \I__10801\ : Odrv4
    port map (
            O => \N__46667\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10800\ : Odrv4
    port map (
            O => \N__46664\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10799\ : Odrv4
    port map (
            O => \N__46661\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10798\ : Odrv12
    port map (
            O => \N__46658\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10797\ : InMux
    port map (
            O => \N__46649\,
            I => \N__46645\
        );

    \I__10796\ : CascadeMux
    port map (
            O => \N__46648\,
            I => \N__46642\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__46645\,
            I => \N__46639\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46635\
        );

    \I__10793\ : Span4Mux_h
    port map (
            O => \N__46639\,
            I => \N__46632\
        );

    \I__10792\ : InMux
    port map (
            O => \N__46638\,
            I => \N__46629\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__46635\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__10790\ : Odrv4
    port map (
            O => \N__46632\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__46629\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46622\,
            I => \N__46619\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__46619\,
            I => \N__46616\
        );

    \I__10786\ : Odrv12
    port map (
            O => \N__46616\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__10785\ : InMux
    port map (
            O => \N__46613\,
            I => \N__46606\
        );

    \I__10784\ : InMux
    port map (
            O => \N__46612\,
            I => \N__46606\
        );

    \I__10783\ : InMux
    port map (
            O => \N__46611\,
            I => \N__46603\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__46606\,
            I => \N__46600\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46603\,
            I => \N__46597\
        );

    \I__10780\ : Span4Mux_h
    port map (
            O => \N__46600\,
            I => \N__46594\
        );

    \I__10779\ : Span4Mux_h
    port map (
            O => \N__46597\,
            I => \N__46588\
        );

    \I__10778\ : Span4Mux_v
    port map (
            O => \N__46594\,
            I => \N__46588\
        );

    \I__10777\ : InMux
    port map (
            O => \N__46593\,
            I => \N__46585\
        );

    \I__10776\ : Odrv4
    port map (
            O => \N__46588\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__46585\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__10774\ : InMux
    port map (
            O => \N__46580\,
            I => \N__46573\
        );

    \I__10773\ : InMux
    port map (
            O => \N__46579\,
            I => \N__46573\
        );

    \I__10772\ : InMux
    port map (
            O => \N__46578\,
            I => \N__46570\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__46573\,
            I => \N__46567\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46570\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__46567\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__10768\ : InMux
    port map (
            O => \N__46562\,
            I => \N__46559\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__46559\,
            I => \N__46556\
        );

    \I__10766\ : Span4Mux_h
    port map (
            O => \N__46556\,
            I => \N__46553\
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__46553\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__10764\ : CascadeMux
    port map (
            O => \N__46550\,
            I => \N__46547\
        );

    \I__10763\ : InMux
    port map (
            O => \N__46547\,
            I => \N__46542\
        );

    \I__10762\ : InMux
    port map (
            O => \N__46546\,
            I => \N__46539\
        );

    \I__10761\ : InMux
    port map (
            O => \N__46545\,
            I => \N__46536\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__46542\,
            I => \N__46533\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46539\,
            I => \N__46530\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__46536\,
            I => \N__46527\
        );

    \I__10757\ : Span4Mux_v
    port map (
            O => \N__46533\,
            I => \N__46522\
        );

    \I__10756\ : Span4Mux_h
    port map (
            O => \N__46530\,
            I => \N__46522\
        );

    \I__10755\ : Span4Mux_v
    port map (
            O => \N__46527\,
            I => \N__46518\
        );

    \I__10754\ : Span4Mux_v
    port map (
            O => \N__46522\,
            I => \N__46515\
        );

    \I__10753\ : InMux
    port map (
            O => \N__46521\,
            I => \N__46512\
        );

    \I__10752\ : Odrv4
    port map (
            O => \N__46518\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10751\ : Odrv4
    port map (
            O => \N__46515\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__46512\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46505\,
            I => \N__46502\
        );

    \I__10748\ : LocalMux
    port map (
            O => \N__46502\,
            I => \N__46497\
        );

    \I__10747\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46494\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46500\,
            I => \N__46491\
        );

    \I__10745\ : Odrv4
    port map (
            O => \N__46497\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__46494\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__46491\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__10742\ : InMux
    port map (
            O => \N__46484\,
            I => \N__46481\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__46481\,
            I => \N__46478\
        );

    \I__10740\ : Odrv4
    port map (
            O => \N__46478\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__10739\ : InMux
    port map (
            O => \N__46475\,
            I => \N__46472\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__46472\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__10737\ : InMux
    port map (
            O => \N__46469\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__10736\ : CascadeMux
    port map (
            O => \N__46466\,
            I => \N__46463\
        );

    \I__10735\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46456\
        );

    \I__10734\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46453\
        );

    \I__10733\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46446\
        );

    \I__10732\ : InMux
    port map (
            O => \N__46460\,
            I => \N__46446\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46459\,
            I => \N__46446\
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__46456\,
            I => \N__46433\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__46453\,
            I => \N__46433\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__46446\,
            I => \N__46430\
        );

    \I__10727\ : InMux
    port map (
            O => \N__46445\,
            I => \N__46413\
        );

    \I__10726\ : InMux
    port map (
            O => \N__46444\,
            I => \N__46413\
        );

    \I__10725\ : InMux
    port map (
            O => \N__46443\,
            I => \N__46413\
        );

    \I__10724\ : InMux
    port map (
            O => \N__46442\,
            I => \N__46413\
        );

    \I__10723\ : InMux
    port map (
            O => \N__46441\,
            I => \N__46413\
        );

    \I__10722\ : InMux
    port map (
            O => \N__46440\,
            I => \N__46413\
        );

    \I__10721\ : InMux
    port map (
            O => \N__46439\,
            I => \N__46413\
        );

    \I__10720\ : InMux
    port map (
            O => \N__46438\,
            I => \N__46413\
        );

    \I__10719\ : Span4Mux_v
    port map (
            O => \N__46433\,
            I => \N__46406\
        );

    \I__10718\ : Span4Mux_v
    port map (
            O => \N__46430\,
            I => \N__46406\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__46413\,
            I => \N__46406\
        );

    \I__10716\ : Odrv4
    port map (
            O => \N__46406\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10715\ : InMux
    port map (
            O => \N__46403\,
            I => \N__46400\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__46400\,
            I => \N__46397\
        );

    \I__10713\ : Odrv12
    port map (
            O => \N__46397\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__10712\ : InMux
    port map (
            O => \N__46394\,
            I => \N__46390\
        );

    \I__10711\ : CascadeMux
    port map (
            O => \N__46393\,
            I => \N__46387\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__46390\,
            I => \N__46384\
        );

    \I__10709\ : InMux
    port map (
            O => \N__46387\,
            I => \N__46381\
        );

    \I__10708\ : Span4Mux_h
    port map (
            O => \N__46384\,
            I => \N__46377\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__46381\,
            I => \N__46374\
        );

    \I__10706\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46371\
        );

    \I__10705\ : Span4Mux_v
    port map (
            O => \N__46377\,
            I => \N__46366\
        );

    \I__10704\ : Span4Mux_h
    port map (
            O => \N__46374\,
            I => \N__46366\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__46371\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10702\ : Odrv4
    port map (
            O => \N__46366\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10701\ : InMux
    port map (
            O => \N__46361\,
            I => \N__46358\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__46358\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__10699\ : CascadeMux
    port map (
            O => \N__46355\,
            I => \N__46350\
        );

    \I__10698\ : CascadeMux
    port map (
            O => \N__46354\,
            I => \N__46346\
        );

    \I__10697\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46341\
        );

    \I__10696\ : InMux
    port map (
            O => \N__46350\,
            I => \N__46341\
        );

    \I__10695\ : CascadeMux
    port map (
            O => \N__46349\,
            I => \N__46338\
        );

    \I__10694\ : InMux
    port map (
            O => \N__46346\,
            I => \N__46335\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__46341\,
            I => \N__46332\
        );

    \I__10692\ : InMux
    port map (
            O => \N__46338\,
            I => \N__46329\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__46335\,
            I => \N__46326\
        );

    \I__10690\ : Odrv12
    port map (
            O => \N__46332\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__46329\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10688\ : Odrv4
    port map (
            O => \N__46326\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10687\ : InMux
    port map (
            O => \N__46319\,
            I => \N__46316\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__46316\,
            I => \N__46313\
        );

    \I__10685\ : Span4Mux_h
    port map (
            O => \N__46313\,
            I => \N__46310\
        );

    \I__10684\ : Odrv4
    port map (
            O => \N__46310\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__10683\ : CascadeMux
    port map (
            O => \N__46307\,
            I => \N__46304\
        );

    \I__10682\ : InMux
    port map (
            O => \N__46304\,
            I => \N__46295\
        );

    \I__10681\ : InMux
    port map (
            O => \N__46303\,
            I => \N__46295\
        );

    \I__10680\ : InMux
    port map (
            O => \N__46302\,
            I => \N__46295\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__46295\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__10678\ : InMux
    port map (
            O => \N__46292\,
            I => \N__46280\
        );

    \I__10677\ : InMux
    port map (
            O => \N__46291\,
            I => \N__46280\
        );

    \I__10676\ : InMux
    port map (
            O => \N__46290\,
            I => \N__46280\
        );

    \I__10675\ : InMux
    port map (
            O => \N__46289\,
            I => \N__46280\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__46280\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__10673\ : InMux
    port map (
            O => \N__46277\,
            I => \N__46274\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__46274\,
            I => \N__46271\
        );

    \I__10671\ : Odrv12
    port map (
            O => \N__46271\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__10670\ : CascadeMux
    port map (
            O => \N__46268\,
            I => \N__46263\
        );

    \I__10669\ : CascadeMux
    port map (
            O => \N__46267\,
            I => \N__46260\
        );

    \I__10668\ : InMux
    port map (
            O => \N__46266\,
            I => \N__46257\
        );

    \I__10667\ : InMux
    port map (
            O => \N__46263\,
            I => \N__46254\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46260\,
            I => \N__46251\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__46257\,
            I => \N__46248\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__46254\,
            I => \N__46245\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__46251\,
            I => \N__46242\
        );

    \I__10662\ : Span4Mux_h
    port map (
            O => \N__46248\,
            I => \N__46239\
        );

    \I__10661\ : Span4Mux_v
    port map (
            O => \N__46245\,
            I => \N__46233\
        );

    \I__10660\ : Span4Mux_v
    port map (
            O => \N__46242\,
            I => \N__46233\
        );

    \I__10659\ : Span4Mux_v
    port map (
            O => \N__46239\,
            I => \N__46230\
        );

    \I__10658\ : InMux
    port map (
            O => \N__46238\,
            I => \N__46227\
        );

    \I__10657\ : Odrv4
    port map (
            O => \N__46233\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10656\ : Odrv4
    port map (
            O => \N__46230\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__46227\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__10654\ : InMux
    port map (
            O => \N__46220\,
            I => \N__46215\
        );

    \I__10653\ : InMux
    port map (
            O => \N__46219\,
            I => \N__46212\
        );

    \I__10652\ : InMux
    port map (
            O => \N__46218\,
            I => \N__46209\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__46215\,
            I => \N__46206\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__46212\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__46209\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__10648\ : Odrv4
    port map (
            O => \N__46206\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__10647\ : InMux
    port map (
            O => \N__46199\,
            I => \N__46196\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__46196\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__10645\ : InMux
    port map (
            O => \N__46193\,
            I => \N__46187\
        );

    \I__10644\ : InMux
    port map (
            O => \N__46192\,
            I => \N__46187\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__46187\,
            I => \N__46184\
        );

    \I__10642\ : Span4Mux_h
    port map (
            O => \N__46184\,
            I => \N__46180\
        );

    \I__10641\ : InMux
    port map (
            O => \N__46183\,
            I => \N__46177\
        );

    \I__10640\ : Odrv4
    port map (
            O => \N__46180\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__46177\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__10638\ : InMux
    port map (
            O => \N__46172\,
            I => \N__46169\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__46169\,
            I => \N__46166\
        );

    \I__10636\ : Span4Mux_v
    port map (
            O => \N__46166\,
            I => \N__46163\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__46163\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__10634\ : CascadeMux
    port map (
            O => \N__46160\,
            I => \N__46157\
        );

    \I__10633\ : InMux
    port map (
            O => \N__46157\,
            I => \N__46154\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__46154\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__46151\,
            I => \N__46142\
        );

    \I__10630\ : CascadeMux
    port map (
            O => \N__46150\,
            I => \N__46139\
        );

    \I__10629\ : CascadeMux
    port map (
            O => \N__46149\,
            I => \N__46136\
        );

    \I__10628\ : CascadeMux
    port map (
            O => \N__46148\,
            I => \N__46133\
        );

    \I__10627\ : CascadeMux
    port map (
            O => \N__46147\,
            I => \N__46130\
        );

    \I__10626\ : CascadeMux
    port map (
            O => \N__46146\,
            I => \N__46126\
        );

    \I__10625\ : CascadeMux
    port map (
            O => \N__46145\,
            I => \N__46123\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46142\,
            I => \N__46104\
        );

    \I__10623\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46104\
        );

    \I__10622\ : InMux
    port map (
            O => \N__46136\,
            I => \N__46104\
        );

    \I__10621\ : InMux
    port map (
            O => \N__46133\,
            I => \N__46104\
        );

    \I__10620\ : InMux
    port map (
            O => \N__46130\,
            I => \N__46095\
        );

    \I__10619\ : InMux
    port map (
            O => \N__46129\,
            I => \N__46095\
        );

    \I__10618\ : InMux
    port map (
            O => \N__46126\,
            I => \N__46095\
        );

    \I__10617\ : InMux
    port map (
            O => \N__46123\,
            I => \N__46095\
        );

    \I__10616\ : CascadeMux
    port map (
            O => \N__46122\,
            I => \N__46091\
        );

    \I__10615\ : CascadeMux
    port map (
            O => \N__46121\,
            I => \N__46088\
        );

    \I__10614\ : CascadeMux
    port map (
            O => \N__46120\,
            I => \N__46085\
        );

    \I__10613\ : CascadeMux
    port map (
            O => \N__46119\,
            I => \N__46082\
        );

    \I__10612\ : CascadeMux
    port map (
            O => \N__46118\,
            I => \N__46078\
        );

    \I__10611\ : CascadeMux
    port map (
            O => \N__46117\,
            I => \N__46075\
        );

    \I__10610\ : CascadeMux
    port map (
            O => \N__46116\,
            I => \N__46072\
        );

    \I__10609\ : CascadeMux
    port map (
            O => \N__46115\,
            I => \N__46069\
        );

    \I__10608\ : CascadeMux
    port map (
            O => \N__46114\,
            I => \N__46065\
        );

    \I__10607\ : CascadeMux
    port map (
            O => \N__46113\,
            I => \N__46062\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__46104\,
            I => \N__46056\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__46095\,
            I => \N__46053\
        );

    \I__10604\ : InMux
    port map (
            O => \N__46094\,
            I => \N__46042\
        );

    \I__10603\ : InMux
    port map (
            O => \N__46091\,
            I => \N__46042\
        );

    \I__10602\ : InMux
    port map (
            O => \N__46088\,
            I => \N__46042\
        );

    \I__10601\ : InMux
    port map (
            O => \N__46085\,
            I => \N__46042\
        );

    \I__10600\ : InMux
    port map (
            O => \N__46082\,
            I => \N__46042\
        );

    \I__10599\ : InMux
    port map (
            O => \N__46081\,
            I => \N__46032\
        );

    \I__10598\ : InMux
    port map (
            O => \N__46078\,
            I => \N__46017\
        );

    \I__10597\ : InMux
    port map (
            O => \N__46075\,
            I => \N__46017\
        );

    \I__10596\ : InMux
    port map (
            O => \N__46072\,
            I => \N__46017\
        );

    \I__10595\ : InMux
    port map (
            O => \N__46069\,
            I => \N__46008\
        );

    \I__10594\ : InMux
    port map (
            O => \N__46068\,
            I => \N__46008\
        );

    \I__10593\ : InMux
    port map (
            O => \N__46065\,
            I => \N__46008\
        );

    \I__10592\ : InMux
    port map (
            O => \N__46062\,
            I => \N__46008\
        );

    \I__10591\ : CascadeMux
    port map (
            O => \N__46061\,
            I => \N__46005\
        );

    \I__10590\ : CascadeMux
    port map (
            O => \N__46060\,
            I => \N__46002\
        );

    \I__10589\ : CascadeMux
    port map (
            O => \N__46059\,
            I => \N__45999\
        );

    \I__10588\ : Span4Mux_v
    port map (
            O => \N__46056\,
            I => \N__45992\
        );

    \I__10587\ : Span4Mux_h
    port map (
            O => \N__46053\,
            I => \N__45992\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__46042\,
            I => \N__45992\
        );

    \I__10585\ : CascadeMux
    port map (
            O => \N__46041\,
            I => \N__45989\
        );

    \I__10584\ : CascadeMux
    port map (
            O => \N__46040\,
            I => \N__45986\
        );

    \I__10583\ : CascadeMux
    port map (
            O => \N__46039\,
            I => \N__45983\
        );

    \I__10582\ : CascadeMux
    port map (
            O => \N__46038\,
            I => \N__45980\
        );

    \I__10581\ : CascadeMux
    port map (
            O => \N__46037\,
            I => \N__45977\
        );

    \I__10580\ : CascadeMux
    port map (
            O => \N__46036\,
            I => \N__45974\
        );

    \I__10579\ : CascadeMux
    port map (
            O => \N__46035\,
            I => \N__45971\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__46032\,
            I => \N__45968\
        );

    \I__10577\ : InMux
    port map (
            O => \N__46031\,
            I => \N__45963\
        );

    \I__10576\ : InMux
    port map (
            O => \N__46030\,
            I => \N__45956\
        );

    \I__10575\ : InMux
    port map (
            O => \N__46029\,
            I => \N__45956\
        );

    \I__10574\ : InMux
    port map (
            O => \N__46028\,
            I => \N__45956\
        );

    \I__10573\ : InMux
    port map (
            O => \N__46027\,
            I => \N__45947\
        );

    \I__10572\ : InMux
    port map (
            O => \N__46026\,
            I => \N__45947\
        );

    \I__10571\ : InMux
    port map (
            O => \N__46025\,
            I => \N__45947\
        );

    \I__10570\ : InMux
    port map (
            O => \N__46024\,
            I => \N__45947\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__46017\,
            I => \N__45942\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__46008\,
            I => \N__45942\
        );

    \I__10567\ : InMux
    port map (
            O => \N__46005\,
            I => \N__45935\
        );

    \I__10566\ : InMux
    port map (
            O => \N__46002\,
            I => \N__45935\
        );

    \I__10565\ : InMux
    port map (
            O => \N__45999\,
            I => \N__45935\
        );

    \I__10564\ : Span4Mux_v
    port map (
            O => \N__45992\,
            I => \N__45932\
        );

    \I__10563\ : InMux
    port map (
            O => \N__45989\,
            I => \N__45925\
        );

    \I__10562\ : InMux
    port map (
            O => \N__45986\,
            I => \N__45925\
        );

    \I__10561\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45925\
        );

    \I__10560\ : InMux
    port map (
            O => \N__45980\,
            I => \N__45916\
        );

    \I__10559\ : InMux
    port map (
            O => \N__45977\,
            I => \N__45916\
        );

    \I__10558\ : InMux
    port map (
            O => \N__45974\,
            I => \N__45916\
        );

    \I__10557\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45916\
        );

    \I__10556\ : Span4Mux_v
    port map (
            O => \N__45968\,
            I => \N__45913\
        );

    \I__10555\ : InMux
    port map (
            O => \N__45967\,
            I => \N__45909\
        );

    \I__10554\ : CascadeMux
    port map (
            O => \N__45966\,
            I => \N__45904\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__45963\,
            I => \N__45897\
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__45956\,
            I => \N__45897\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__45947\,
            I => \N__45897\
        );

    \I__10550\ : Span4Mux_v
    port map (
            O => \N__45942\,
            I => \N__45878\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__45935\,
            I => \N__45878\
        );

    \I__10548\ : Span4Mux_v
    port map (
            O => \N__45932\,
            I => \N__45878\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__45925\,
            I => \N__45878\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__45916\,
            I => \N__45878\
        );

    \I__10545\ : Span4Mux_h
    port map (
            O => \N__45913\,
            I => \N__45875\
        );

    \I__10544\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45872\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__45909\,
            I => \N__45869\
        );

    \I__10542\ : InMux
    port map (
            O => \N__45908\,
            I => \N__45866\
        );

    \I__10541\ : InMux
    port map (
            O => \N__45907\,
            I => \N__45861\
        );

    \I__10540\ : InMux
    port map (
            O => \N__45904\,
            I => \N__45861\
        );

    \I__10539\ : Span4Mux_v
    port map (
            O => \N__45897\,
            I => \N__45858\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45896\,
            I => \N__45849\
        );

    \I__10537\ : InMux
    port map (
            O => \N__45895\,
            I => \N__45849\
        );

    \I__10536\ : InMux
    port map (
            O => \N__45894\,
            I => \N__45849\
        );

    \I__10535\ : InMux
    port map (
            O => \N__45893\,
            I => \N__45840\
        );

    \I__10534\ : InMux
    port map (
            O => \N__45892\,
            I => \N__45840\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45891\,
            I => \N__45840\
        );

    \I__10532\ : InMux
    port map (
            O => \N__45890\,
            I => \N__45840\
        );

    \I__10531\ : CascadeMux
    port map (
            O => \N__45889\,
            I => \N__45837\
        );

    \I__10530\ : Sp12to4
    port map (
            O => \N__45878\,
            I => \N__45833\
        );

    \I__10529\ : Span4Mux_v
    port map (
            O => \N__45875\,
            I => \N__45830\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__45872\,
            I => \N__45825\
        );

    \I__10527\ : Span4Mux_s1_v
    port map (
            O => \N__45869\,
            I => \N__45825\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__45866\,
            I => \N__45822\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__45861\,
            I => \N__45819\
        );

    \I__10524\ : Span4Mux_v
    port map (
            O => \N__45858\,
            I => \N__45816\
        );

    \I__10523\ : InMux
    port map (
            O => \N__45857\,
            I => \N__45813\
        );

    \I__10522\ : CascadeMux
    port map (
            O => \N__45856\,
            I => \N__45810\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__45849\,
            I => \N__45805\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__45840\,
            I => \N__45805\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45837\,
            I => \N__45800\
        );

    \I__10518\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45800\
        );

    \I__10517\ : Span12Mux_v
    port map (
            O => \N__45833\,
            I => \N__45795\
        );

    \I__10516\ : Sp12to4
    port map (
            O => \N__45830\,
            I => \N__45795\
        );

    \I__10515\ : Span4Mux_v
    port map (
            O => \N__45825\,
            I => \N__45790\
        );

    \I__10514\ : Span4Mux_v
    port map (
            O => \N__45822\,
            I => \N__45790\
        );

    \I__10513\ : Span12Mux_v
    port map (
            O => \N__45819\,
            I => \N__45787\
        );

    \I__10512\ : Sp12to4
    port map (
            O => \N__45816\,
            I => \N__45782\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__45813\,
            I => \N__45782\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45810\,
            I => \N__45779\
        );

    \I__10509\ : Span4Mux_s2_h
    port map (
            O => \N__45805\,
            I => \N__45774\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__45800\,
            I => \N__45774\
        );

    \I__10507\ : Span12Mux_h
    port map (
            O => \N__45795\,
            I => \N__45771\
        );

    \I__10506\ : Span4Mux_v
    port map (
            O => \N__45790\,
            I => \N__45768\
        );

    \I__10505\ : Span12Mux_h
    port map (
            O => \N__45787\,
            I => \N__45759\
        );

    \I__10504\ : Span12Mux_s2_h
    port map (
            O => \N__45782\,
            I => \N__45759\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__45779\,
            I => \N__45759\
        );

    \I__10502\ : Sp12to4
    port map (
            O => \N__45774\,
            I => \N__45759\
        );

    \I__10501\ : Odrv12
    port map (
            O => \N__45771\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10500\ : Odrv4
    port map (
            O => \N__45768\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10499\ : Odrv12
    port map (
            O => \N__45759\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10498\ : CascadeMux
    port map (
            O => \N__45752\,
            I => \N__45749\
        );

    \I__10497\ : InMux
    port map (
            O => \N__45749\,
            I => \N__45746\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__45746\,
            I => \N__45743\
        );

    \I__10495\ : Odrv4
    port map (
            O => \N__45743\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__10494\ : InMux
    port map (
            O => \N__45740\,
            I => \N__45737\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__45737\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45734\,
            I => \N__45731\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__45731\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__10490\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45725\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__45725\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45722\,
            I => \N__45719\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__45719\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__10486\ : InMux
    port map (
            O => \N__45716\,
            I => \N__45713\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45713\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__10484\ : InMux
    port map (
            O => \N__45710\,
            I => \N__45707\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__45707\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__10482\ : CascadeMux
    port map (
            O => \N__45704\,
            I => \N__45701\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45701\,
            I => \N__45698\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__45698\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45692\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__45692\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45689\,
            I => \N__45686\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__45686\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45683\,
            I => \N__45680\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__45680\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__10473\ : InMux
    port map (
            O => \N__45677\,
            I => \N__45674\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__45674\,
            I => \N__45671\
        );

    \I__10471\ : Odrv12
    port map (
            O => \N__45671\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45663\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45667\,
            I => \N__45660\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45666\,
            I => \N__45657\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__45663\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__45660\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__45657\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10464\ : CascadeMux
    port map (
            O => \N__45650\,
            I => \N__45646\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45649\,
            I => \N__45643\
        );

    \I__10462\ : InMux
    port map (
            O => \N__45646\,
            I => \N__45640\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__45643\,
            I => \N__45637\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__45640\,
            I => \N__45634\
        );

    \I__10459\ : Span4Mux_h
    port map (
            O => \N__45637\,
            I => \N__45631\
        );

    \I__10458\ : Span4Mux_v
    port map (
            O => \N__45634\,
            I => \N__45628\
        );

    \I__10457\ : Span4Mux_h
    port map (
            O => \N__45631\,
            I => \N__45625\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__45628\,
            I => \N__45622\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__45625\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__10454\ : Odrv4
    port map (
            O => \N__45622\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45617\,
            I => \N__45612\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45609\
        );

    \I__10451\ : InMux
    port map (
            O => \N__45615\,
            I => \N__45606\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__45612\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45609\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__45606\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10447\ : InMux
    port map (
            O => \N__45599\,
            I => \N__45596\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45596\,
            I => \N__45591\
        );

    \I__10445\ : InMux
    port map (
            O => \N__45595\,
            I => \N__45588\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45594\,
            I => \N__45585\
        );

    \I__10443\ : Span4Mux_h
    port map (
            O => \N__45591\,
            I => \N__45580\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__45588\,
            I => \N__45580\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__45585\,
            I => \N__45577\
        );

    \I__10440\ : Span4Mux_h
    port map (
            O => \N__45580\,
            I => \N__45574\
        );

    \I__10439\ : Odrv12
    port map (
            O => \N__45577\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__10438\ : Odrv4
    port map (
            O => \N__45574\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__10437\ : CEMux
    port map (
            O => \N__45569\,
            I => \N__45551\
        );

    \I__10436\ : CEMux
    port map (
            O => \N__45568\,
            I => \N__45551\
        );

    \I__10435\ : CEMux
    port map (
            O => \N__45567\,
            I => \N__45551\
        );

    \I__10434\ : CEMux
    port map (
            O => \N__45566\,
            I => \N__45551\
        );

    \I__10433\ : CEMux
    port map (
            O => \N__45565\,
            I => \N__45551\
        );

    \I__10432\ : CEMux
    port map (
            O => \N__45564\,
            I => \N__45551\
        );

    \I__10431\ : GlobalMux
    port map (
            O => \N__45551\,
            I => \N__45548\
        );

    \I__10430\ : gio2CtrlBuf
    port map (
            O => \N__45548\,
            I => \delay_measurement_inst.delay_tr_timer.N_304_i_g\
        );

    \I__10429\ : InMux
    port map (
            O => \N__45545\,
            I => \N__45542\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45542\,
            I => \N__45538\
        );

    \I__10427\ : InMux
    port map (
            O => \N__45541\,
            I => \N__45535\
        );

    \I__10426\ : Span4Mux_s1_v
    port map (
            O => \N__45538\,
            I => \N__45530\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__45535\,
            I => \N__45530\
        );

    \I__10424\ : Span4Mux_v
    port map (
            O => \N__45530\,
            I => \N__45527\
        );

    \I__10423\ : Span4Mux_h
    port map (
            O => \N__45527\,
            I => \N__45524\
        );

    \I__10422\ : Sp12to4
    port map (
            O => \N__45524\,
            I => \N__45520\
        );

    \I__10421\ : InMux
    port map (
            O => \N__45523\,
            I => \N__45517\
        );

    \I__10420\ : Span12Mux_v
    port map (
            O => \N__45520\,
            I => \N__45514\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__45517\,
            I => \N__45511\
        );

    \I__10418\ : Span12Mux_v
    port map (
            O => \N__45514\,
            I => \N__45507\
        );

    \I__10417\ : Span12Mux_h
    port map (
            O => \N__45511\,
            I => \N__45504\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45501\
        );

    \I__10415\ : Span12Mux_h
    port map (
            O => \N__45507\,
            I => \N__45496\
        );

    \I__10414\ : Span12Mux_v
    port map (
            O => \N__45504\,
            I => \N__45496\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__45501\,
            I => \N__45493\
        );

    \I__10412\ : Odrv12
    port map (
            O => \N__45496\,
            I => start_stop_c
        );

    \I__10411\ : Odrv12
    port map (
            O => \N__45493\,
            I => start_stop_c
        );

    \I__10410\ : InMux
    port map (
            O => \N__45488\,
            I => \N__45483\
        );

    \I__10409\ : InMux
    port map (
            O => \N__45487\,
            I => \N__45476\
        );

    \I__10408\ : InMux
    port map (
            O => \N__45486\,
            I => \N__45476\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__45483\,
            I => \N__45473\
        );

    \I__10406\ : InMux
    port map (
            O => \N__45482\,
            I => \N__45470\
        );

    \I__10405\ : InMux
    port map (
            O => \N__45481\,
            I => \N__45467\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__45476\,
            I => \N__45464\
        );

    \I__10403\ : Span4Mux_v
    port map (
            O => \N__45473\,
            I => \N__45459\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__45470\,
            I => \N__45459\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__45467\,
            I => \N__45455\
        );

    \I__10400\ : Span4Mux_h
    port map (
            O => \N__45464\,
            I => \N__45452\
        );

    \I__10399\ : Span4Mux_v
    port map (
            O => \N__45459\,
            I => \N__45449\
        );

    \I__10398\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45446\
        );

    \I__10397\ : Span4Mux_v
    port map (
            O => \N__45455\,
            I => \N__45439\
        );

    \I__10396\ : Span4Mux_v
    port map (
            O => \N__45452\,
            I => \N__45439\
        );

    \I__10395\ : Span4Mux_h
    port map (
            O => \N__45449\,
            I => \N__45439\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__45446\,
            I => phase_controller_inst1_state_4
        );

    \I__10393\ : Odrv4
    port map (
            O => \N__45439\,
            I => phase_controller_inst1_state_4
        );

    \I__10392\ : InMux
    port map (
            O => \N__45434\,
            I => \N__45430\
        );

    \I__10391\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45427\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__45430\,
            I => \N__45424\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__45427\,
            I => \N__45421\
        );

    \I__10388\ : Span4Mux_v
    port map (
            O => \N__45424\,
            I => \N__45418\
        );

    \I__10387\ : Span4Mux_h
    port map (
            O => \N__45421\,
            I => \N__45415\
        );

    \I__10386\ : Span4Mux_v
    port map (
            O => \N__45418\,
            I => \N__45412\
        );

    \I__10385\ : Span4Mux_v
    port map (
            O => \N__45415\,
            I => \N__45409\
        );

    \I__10384\ : Odrv4
    port map (
            O => \N__45412\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__10383\ : Odrv4
    port map (
            O => \N__45409\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__10382\ : CascadeMux
    port map (
            O => \N__45404\,
            I => \N__45401\
        );

    \I__10381\ : InMux
    port map (
            O => \N__45401\,
            I => \N__45398\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__45398\,
            I => \N__45393\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45397\,
            I => \N__45388\
        );

    \I__10378\ : InMux
    port map (
            O => \N__45396\,
            I => \N__45388\
        );

    \I__10377\ : Span4Mux_v
    port map (
            O => \N__45393\,
            I => \N__45385\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__45388\,
            I => \N__45382\
        );

    \I__10375\ : Odrv4
    port map (
            O => \N__45385\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__45382\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__10373\ : InMux
    port map (
            O => \N__45377\,
            I => \N__45374\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__45374\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__10371\ : InMux
    port map (
            O => \N__45371\,
            I => \N__45368\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__45368\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__10369\ : InMux
    port map (
            O => \N__45365\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__10368\ : InMux
    port map (
            O => \N__45362\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__10367\ : CascadeMux
    port map (
            O => \N__45359\,
            I => \N__45356\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45356\,
            I => \N__45353\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__45353\,
            I => \N__45350\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__45350\,
            I => \N__45347\
        );

    \I__10363\ : Span4Mux_v
    port map (
            O => \N__45347\,
            I => \N__45344\
        );

    \I__10362\ : Odrv4
    port map (
            O => \N__45344\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__10361\ : CascadeMux
    port map (
            O => \N__45341\,
            I => \N__45338\
        );

    \I__10360\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45335\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__45335\,
            I => \N__45332\
        );

    \I__10358\ : Span4Mux_h
    port map (
            O => \N__45332\,
            I => \N__45329\
        );

    \I__10357\ : Odrv4
    port map (
            O => \N__45329\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__10356\ : CascadeMux
    port map (
            O => \N__45326\,
            I => \N__45321\
        );

    \I__10355\ : InMux
    port map (
            O => \N__45325\,
            I => \N__45318\
        );

    \I__10354\ : InMux
    port map (
            O => \N__45324\,
            I => \N__45315\
        );

    \I__10353\ : InMux
    port map (
            O => \N__45321\,
            I => \N__45312\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__45318\,
            I => \N__45309\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__45315\,
            I => \N__45306\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__45312\,
            I => \N__45303\
        );

    \I__10349\ : Span4Mux_h
    port map (
            O => \N__45309\,
            I => \N__45300\
        );

    \I__10348\ : Span4Mux_h
    port map (
            O => \N__45306\,
            I => \N__45295\
        );

    \I__10347\ : Span4Mux_h
    port map (
            O => \N__45303\,
            I => \N__45295\
        );

    \I__10346\ : Odrv4
    port map (
            O => \N__45300\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10345\ : Odrv4
    port map (
            O => \N__45295\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10344\ : CascadeMux
    port map (
            O => \N__45290\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__10343\ : CascadeMux
    port map (
            O => \N__45287\,
            I => \N__45284\
        );

    \I__10342\ : InMux
    port map (
            O => \N__45284\,
            I => \N__45278\
        );

    \I__10341\ : InMux
    port map (
            O => \N__45283\,
            I => \N__45273\
        );

    \I__10340\ : InMux
    port map (
            O => \N__45282\,
            I => \N__45273\
        );

    \I__10339\ : InMux
    port map (
            O => \N__45281\,
            I => \N__45270\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__45278\,
            I => \N__45267\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__45273\,
            I => \N__45264\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__45270\,
            I => \N__45261\
        );

    \I__10335\ : Span4Mux_v
    port map (
            O => \N__45267\,
            I => \N__45258\
        );

    \I__10334\ : Span12Mux_s10_h
    port map (
            O => \N__45264\,
            I => \N__45255\
        );

    \I__10333\ : Span4Mux_h
    port map (
            O => \N__45261\,
            I => \N__45252\
        );

    \I__10332\ : Odrv4
    port map (
            O => \N__45258\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10331\ : Odrv12
    port map (
            O => \N__45255\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10330\ : Odrv4
    port map (
            O => \N__45252\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10329\ : InMux
    port map (
            O => \N__45245\,
            I => \N__45242\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__45242\,
            I => \N__45239\
        );

    \I__10327\ : Odrv4
    port map (
            O => \N__45239\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__10326\ : InMux
    port map (
            O => \N__45236\,
            I => \N__45233\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__45233\,
            I => \N__45228\
        );

    \I__10324\ : InMux
    port map (
            O => \N__45232\,
            I => \N__45222\
        );

    \I__10323\ : InMux
    port map (
            O => \N__45231\,
            I => \N__45222\
        );

    \I__10322\ : Span4Mux_v
    port map (
            O => \N__45228\,
            I => \N__45219\
        );

    \I__10321\ : InMux
    port map (
            O => \N__45227\,
            I => \N__45216\
        );

    \I__10320\ : LocalMux
    port map (
            O => \N__45222\,
            I => \N__45213\
        );

    \I__10319\ : Span4Mux_v
    port map (
            O => \N__45219\,
            I => \N__45210\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__45216\,
            I => \N__45207\
        );

    \I__10317\ : Odrv12
    port map (
            O => \N__45213\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10316\ : Odrv4
    port map (
            O => \N__45210\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10315\ : Odrv4
    port map (
            O => \N__45207\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10314\ : InMux
    port map (
            O => \N__45200\,
            I => \N__45197\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__45197\,
            I => \N__45194\
        );

    \I__10312\ : Odrv12
    port map (
            O => \N__45194\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__10311\ : CascadeMux
    port map (
            O => \N__45191\,
            I => \N__45186\
        );

    \I__10310\ : InMux
    port map (
            O => \N__45190\,
            I => \N__45183\
        );

    \I__10309\ : InMux
    port map (
            O => \N__45189\,
            I => \N__45180\
        );

    \I__10308\ : InMux
    port map (
            O => \N__45186\,
            I => \N__45177\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__45183\,
            I => \N__45172\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__45180\,
            I => \N__45172\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__45177\,
            I => \N__45168\
        );

    \I__10304\ : Span4Mux_v
    port map (
            O => \N__45172\,
            I => \N__45165\
        );

    \I__10303\ : InMux
    port map (
            O => \N__45171\,
            I => \N__45162\
        );

    \I__10302\ : Span4Mux_h
    port map (
            O => \N__45168\,
            I => \N__45159\
        );

    \I__10301\ : Span4Mux_v
    port map (
            O => \N__45165\,
            I => \N__45154\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45154\
        );

    \I__10299\ : Odrv4
    port map (
            O => \N__45159\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10298\ : Odrv4
    port map (
            O => \N__45154\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45149\,
            I => \N__45146\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__45146\,
            I => \N__45143\
        );

    \I__10295\ : Odrv12
    port map (
            O => \N__45143\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__10294\ : InMux
    port map (
            O => \N__45140\,
            I => \N__45137\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__45137\,
            I => \N__45134\
        );

    \I__10292\ : Odrv4
    port map (
            O => \N__45134\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__10291\ : InMux
    port map (
            O => \N__45131\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__10290\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45125\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__45125\,
            I => \N__45122\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__45122\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__10287\ : InMux
    port map (
            O => \N__45119\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__10286\ : InMux
    port map (
            O => \N__45116\,
            I => \N__45109\
        );

    \I__10285\ : InMux
    port map (
            O => \N__45115\,
            I => \N__45109\
        );

    \I__10284\ : InMux
    port map (
            O => \N__45114\,
            I => \N__45106\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__45109\,
            I => \N__45103\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__45106\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10281\ : Odrv12
    port map (
            O => \N__45103\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10280\ : InMux
    port map (
            O => \N__45098\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__10279\ : InMux
    port map (
            O => \N__45095\,
            I => \N__45092\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45092\,
            I => \N__45089\
        );

    \I__10277\ : Span4Mux_v
    port map (
            O => \N__45089\,
            I => \N__45086\
        );

    \I__10276\ : Odrv4
    port map (
            O => \N__45086\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__10275\ : InMux
    port map (
            O => \N__45083\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__10274\ : InMux
    port map (
            O => \N__45080\,
            I => \N__45077\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__45077\,
            I => \N__45074\
        );

    \I__10272\ : Odrv4
    port map (
            O => \N__45074\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__10271\ : InMux
    port map (
            O => \N__45071\,
            I => \bfn_17_20_0_\
        );

    \I__10270\ : InMux
    port map (
            O => \N__45068\,
            I => \N__45065\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__45065\,
            I => \N__45062\
        );

    \I__10268\ : Odrv4
    port map (
            O => \N__45062\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__10267\ : InMux
    port map (
            O => \N__45059\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__10266\ : InMux
    port map (
            O => \N__45056\,
            I => \N__45053\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__45053\,
            I => \N__45050\
        );

    \I__10264\ : Span4Mux_h
    port map (
            O => \N__45050\,
            I => \N__45047\
        );

    \I__10263\ : Odrv4
    port map (
            O => \N__45047\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__10262\ : InMux
    port map (
            O => \N__45044\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__10261\ : InMux
    port map (
            O => \N__45041\,
            I => \N__45038\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__45038\,
            I => \N__45035\
        );

    \I__10259\ : Odrv4
    port map (
            O => \N__45035\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__10258\ : InMux
    port map (
            O => \N__45032\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__10257\ : InMux
    port map (
            O => \N__45029\,
            I => \N__45026\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__45026\,
            I => \N__45023\
        );

    \I__10255\ : Odrv4
    port map (
            O => \N__45023\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__10254\ : InMux
    port map (
            O => \N__45020\,
            I => \N__45015\
        );

    \I__10253\ : InMux
    port map (
            O => \N__45019\,
            I => \N__45010\
        );

    \I__10252\ : InMux
    port map (
            O => \N__45018\,
            I => \N__45010\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__45015\,
            I => \N__45007\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__45010\,
            I => \N__45004\
        );

    \I__10249\ : Span4Mux_v
    port map (
            O => \N__45007\,
            I => \N__45001\
        );

    \I__10248\ : Span4Mux_h
    port map (
            O => \N__45004\,
            I => \N__44998\
        );

    \I__10247\ : Odrv4
    port map (
            O => \N__45001\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10246\ : Odrv4
    port map (
            O => \N__44998\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10245\ : InMux
    port map (
            O => \N__44993\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__10244\ : InMux
    port map (
            O => \N__44990\,
            I => \N__44987\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__44987\,
            I => \N__44984\
        );

    \I__10242\ : Span4Mux_h
    port map (
            O => \N__44984\,
            I => \N__44981\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__44981\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__10240\ : InMux
    port map (
            O => \N__44978\,
            I => \N__44971\
        );

    \I__10239\ : InMux
    port map (
            O => \N__44977\,
            I => \N__44971\
        );

    \I__10238\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44968\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__44971\,
            I => \N__44965\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__44968\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10235\ : Odrv4
    port map (
            O => \N__44965\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10234\ : InMux
    port map (
            O => \N__44960\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__10233\ : CascadeMux
    port map (
            O => \N__44957\,
            I => \N__44953\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44956\,
            I => \N__44950\
        );

    \I__10231\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44947\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__44950\,
            I => \N__44944\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__44947\,
            I => \N__44940\
        );

    \I__10228\ : Span4Mux_h
    port map (
            O => \N__44944\,
            I => \N__44937\
        );

    \I__10227\ : InMux
    port map (
            O => \N__44943\,
            I => \N__44934\
        );

    \I__10226\ : Span4Mux_h
    port map (
            O => \N__44940\,
            I => \N__44931\
        );

    \I__10225\ : Span4Mux_v
    port map (
            O => \N__44937\,
            I => \N__44928\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__44934\,
            I => \N__44925\
        );

    \I__10223\ : Odrv4
    port map (
            O => \N__44931\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__10222\ : Odrv4
    port map (
            O => \N__44928\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__10221\ : Odrv12
    port map (
            O => \N__44925\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__10220\ : InMux
    port map (
            O => \N__44918\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__10219\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44912\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__44912\,
            I => \N__44909\
        );

    \I__10217\ : Span4Mux_v
    port map (
            O => \N__44909\,
            I => \N__44906\
        );

    \I__10216\ : Odrv4
    port map (
            O => \N__44906\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__10215\ : CascadeMux
    port map (
            O => \N__44903\,
            I => \N__44899\
        );

    \I__10214\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44893\
        );

    \I__10213\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44893\
        );

    \I__10212\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44890\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__44893\,
            I => \N__44887\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__44890\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10209\ : Odrv4
    port map (
            O => \N__44887\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10208\ : InMux
    port map (
            O => \N__44882\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44879\,
            I => \N__44876\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__44876\,
            I => \N__44873\
        );

    \I__10205\ : Odrv4
    port map (
            O => \N__44873\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44870\,
            I => \bfn_17_19_0_\
        );

    \I__10203\ : InMux
    port map (
            O => \N__44867\,
            I => \N__44864\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__44864\,
            I => \N__44861\
        );

    \I__10201\ : Span4Mux_v
    port map (
            O => \N__44861\,
            I => \N__44858\
        );

    \I__10200\ : Odrv4
    port map (
            O => \N__44858\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__10199\ : InMux
    port map (
            O => \N__44855\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44852\,
            I => \N__44849\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__44849\,
            I => \N__44846\
        );

    \I__10196\ : Span4Mux_h
    port map (
            O => \N__44846\,
            I => \N__44843\
        );

    \I__10195\ : Span4Mux_v
    port map (
            O => \N__44843\,
            I => \N__44840\
        );

    \I__10194\ : Odrv4
    port map (
            O => \N__44840\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__10193\ : InMux
    port map (
            O => \N__44837\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__10192\ : InMux
    port map (
            O => \N__44834\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__10191\ : InMux
    port map (
            O => \N__44831\,
            I => \N__44828\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__44828\,
            I => \N__44825\
        );

    \I__10189\ : Odrv4
    port map (
            O => \N__44825\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__10188\ : InMux
    port map (
            O => \N__44822\,
            I => \N__44818\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44821\,
            I => \N__44814\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__44818\,
            I => \N__44811\
        );

    \I__10185\ : InMux
    port map (
            O => \N__44817\,
            I => \N__44808\
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__44814\,
            I => \N__44805\
        );

    \I__10183\ : Odrv4
    port map (
            O => \N__44811\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__44808\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__10181\ : Odrv12
    port map (
            O => \N__44805\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__10180\ : InMux
    port map (
            O => \N__44798\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44795\,
            I => \N__44789\
        );

    \I__10178\ : InMux
    port map (
            O => \N__44794\,
            I => \N__44789\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__44789\,
            I => \N__44785\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44788\,
            I => \N__44782\
        );

    \I__10175\ : Span4Mux_v
    port map (
            O => \N__44785\,
            I => \N__44779\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__44782\,
            I => \N__44776\
        );

    \I__10173\ : Odrv4
    port map (
            O => \N__44779\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__10172\ : Odrv4
    port map (
            O => \N__44776\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__10171\ : InMux
    port map (
            O => \N__44771\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__10170\ : InMux
    port map (
            O => \N__44768\,
            I => \N__44765\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__44765\,
            I => \N__44762\
        );

    \I__10168\ : Odrv4
    port map (
            O => \N__44762\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44759\,
            I => \N__44752\
        );

    \I__10166\ : InMux
    port map (
            O => \N__44758\,
            I => \N__44752\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44757\,
            I => \N__44749\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__44752\,
            I => \N__44746\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__44749\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__10162\ : Odrv12
    port map (
            O => \N__44746\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__10161\ : InMux
    port map (
            O => \N__44741\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__10160\ : InMux
    port map (
            O => \N__44738\,
            I => \N__44733\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44737\,
            I => \N__44730\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44736\,
            I => \N__44727\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__44733\,
            I => \N__44724\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44730\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__44727\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__10154\ : Odrv4
    port map (
            O => \N__44724\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__10153\ : InMux
    port map (
            O => \N__44717\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__10152\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44711\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__44711\,
            I => \N__44708\
        );

    \I__10150\ : Odrv4
    port map (
            O => \N__44708\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44705\,
            I => \N__44698\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44704\,
            I => \N__44698\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44703\,
            I => \N__44695\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__44698\,
            I => \N__44692\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__44695\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__10144\ : Odrv4
    port map (
            O => \N__44692\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__10143\ : InMux
    port map (
            O => \N__44687\,
            I => \bfn_17_18_0_\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44684\,
            I => \N__44681\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__44681\,
            I => \N__44678\
        );

    \I__10140\ : Odrv4
    port map (
            O => \N__44678\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__10139\ : CascadeMux
    port map (
            O => \N__44675\,
            I => \N__44672\
        );

    \I__10138\ : InMux
    port map (
            O => \N__44672\,
            I => \N__44668\
        );

    \I__10137\ : InMux
    port map (
            O => \N__44671\,
            I => \N__44665\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__44668\,
            I => \N__44661\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__44665\,
            I => \N__44658\
        );

    \I__10134\ : InMux
    port map (
            O => \N__44664\,
            I => \N__44655\
        );

    \I__10133\ : Span4Mux_h
    port map (
            O => \N__44661\,
            I => \N__44652\
        );

    \I__10132\ : Span4Mux_h
    port map (
            O => \N__44658\,
            I => \N__44647\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__44655\,
            I => \N__44647\
        );

    \I__10130\ : Odrv4
    port map (
            O => \N__44652\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10129\ : Odrv4
    port map (
            O => \N__44647\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44642\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__10127\ : InMux
    port map (
            O => \N__44639\,
            I => \N__44636\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__44636\,
            I => \N__44633\
        );

    \I__10125\ : Span4Mux_h
    port map (
            O => \N__44633\,
            I => \N__44630\
        );

    \I__10124\ : Odrv4
    port map (
            O => \N__44630\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44627\,
            I => \N__44623\
        );

    \I__10122\ : InMux
    port map (
            O => \N__44626\,
            I => \N__44619\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__44623\,
            I => \N__44616\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44622\,
            I => \N__44613\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__44619\,
            I => \N__44606\
        );

    \I__10118\ : Span4Mux_h
    port map (
            O => \N__44616\,
            I => \N__44606\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__44613\,
            I => \N__44606\
        );

    \I__10116\ : Odrv4
    port map (
            O => \N__44606\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10115\ : InMux
    port map (
            O => \N__44603\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__10114\ : InMux
    port map (
            O => \N__44600\,
            I => \N__44597\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__44597\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__10112\ : InMux
    port map (
            O => \N__44594\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__10111\ : CascadeMux
    port map (
            O => \N__44591\,
            I => \N__44588\
        );

    \I__10110\ : InMux
    port map (
            O => \N__44588\,
            I => \N__44585\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44585\,
            I => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\
        );

    \I__10108\ : InMux
    port map (
            O => \N__44582\,
            I => \N__44579\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__44579\,
            I => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\
        );

    \I__10106\ : CascadeMux
    port map (
            O => \N__44576\,
            I => \N__44573\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44573\,
            I => \N__44568\
        );

    \I__10104\ : InMux
    port map (
            O => \N__44572\,
            I => \N__44563\
        );

    \I__10103\ : InMux
    port map (
            O => \N__44571\,
            I => \N__44563\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44568\,
            I => \N__44560\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__44563\,
            I => \N__44557\
        );

    \I__10100\ : Span4Mux_h
    port map (
            O => \N__44560\,
            I => \N__44553\
        );

    \I__10099\ : Span12Mux_s10_h
    port map (
            O => \N__44557\,
            I => \N__44550\
        );

    \I__10098\ : InMux
    port map (
            O => \N__44556\,
            I => \N__44547\
        );

    \I__10097\ : Odrv4
    port map (
            O => \N__44553\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10096\ : Odrv12
    port map (
            O => \N__44550\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__44547\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10094\ : CascadeMux
    port map (
            O => \N__44540\,
            I => \N__44537\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44537\,
            I => \N__44532\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44536\,
            I => \N__44529\
        );

    \I__10091\ : InMux
    port map (
            O => \N__44535\,
            I => \N__44526\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__44532\,
            I => \N__44523\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44529\,
            I => \N__44520\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__44526\,
            I => \N__44517\
        );

    \I__10087\ : Span4Mux_h
    port map (
            O => \N__44523\,
            I => \N__44514\
        );

    \I__10086\ : Span4Mux_h
    port map (
            O => \N__44520\,
            I => \N__44511\
        );

    \I__10085\ : Span4Mux_h
    port map (
            O => \N__44517\,
            I => \N__44508\
        );

    \I__10084\ : Span4Mux_v
    port map (
            O => \N__44514\,
            I => \N__44504\
        );

    \I__10083\ : Span4Mux_v
    port map (
            O => \N__44511\,
            I => \N__44501\
        );

    \I__10082\ : Span4Mux_v
    port map (
            O => \N__44508\,
            I => \N__44498\
        );

    \I__10081\ : InMux
    port map (
            O => \N__44507\,
            I => \N__44495\
        );

    \I__10080\ : Odrv4
    port map (
            O => \N__44504\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10079\ : Odrv4
    port map (
            O => \N__44501\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10078\ : Odrv4
    port map (
            O => \N__44498\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__44495\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10076\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44483\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__44483\,
            I => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44480\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__10073\ : InMux
    port map (
            O => \N__44477\,
            I => \N__44474\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__44474\,
            I => \N__44471\
        );

    \I__10071\ : Span4Mux_h
    port map (
            O => \N__44471\,
            I => \N__44468\
        );

    \I__10070\ : Odrv4
    port map (
            O => \N__44468\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44465\,
            I => \N__44462\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__44462\,
            I => \N__44457\
        );

    \I__10067\ : InMux
    port map (
            O => \N__44461\,
            I => \N__44452\
        );

    \I__10066\ : InMux
    port map (
            O => \N__44460\,
            I => \N__44452\
        );

    \I__10065\ : Span4Mux_v
    port map (
            O => \N__44457\,
            I => \N__44449\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__44452\,
            I => \N__44446\
        );

    \I__10063\ : Odrv4
    port map (
            O => \N__44449\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__10062\ : Odrv4
    port map (
            O => \N__44446\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__10061\ : InMux
    port map (
            O => \N__44441\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__10060\ : InMux
    port map (
            O => \N__44438\,
            I => \N__44435\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__44435\,
            I => \N__44432\
        );

    \I__10058\ : Span4Mux_h
    port map (
            O => \N__44432\,
            I => \N__44429\
        );

    \I__10057\ : Odrv4
    port map (
            O => \N__44429\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__10056\ : InMux
    port map (
            O => \N__44426\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__10055\ : InMux
    port map (
            O => \N__44423\,
            I => \N__44420\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__44420\,
            I => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\
        );

    \I__10053\ : InMux
    port map (
            O => \N__44417\,
            I => \N__44413\
        );

    \I__10052\ : InMux
    port map (
            O => \N__44416\,
            I => \N__44409\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__44413\,
            I => \N__44406\
        );

    \I__10050\ : InMux
    port map (
            O => \N__44412\,
            I => \N__44403\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__44409\,
            I => \N__44400\
        );

    \I__10048\ : Span4Mux_h
    port map (
            O => \N__44406\,
            I => \N__44397\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__44403\,
            I => \N__44393\
        );

    \I__10046\ : Span4Mux_h
    port map (
            O => \N__44400\,
            I => \N__44388\
        );

    \I__10045\ : Span4Mux_v
    port map (
            O => \N__44397\,
            I => \N__44388\
        );

    \I__10044\ : InMux
    port map (
            O => \N__44396\,
            I => \N__44385\
        );

    \I__10043\ : Odrv12
    port map (
            O => \N__44393\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10042\ : Odrv4
    port map (
            O => \N__44388\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__44385\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10040\ : CascadeMux
    port map (
            O => \N__44378\,
            I => \N__44373\
        );

    \I__10039\ : InMux
    port map (
            O => \N__44377\,
            I => \N__44368\
        );

    \I__10038\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44368\
        );

    \I__10037\ : InMux
    port map (
            O => \N__44373\,
            I => \N__44365\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__44368\,
            I => \N__44362\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__44365\,
            I => \N__44359\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__44362\,
            I => \N__44356\
        );

    \I__10033\ : Span4Mux_h
    port map (
            O => \N__44359\,
            I => \N__44352\
        );

    \I__10032\ : Span4Mux_v
    port map (
            O => \N__44356\,
            I => \N__44349\
        );

    \I__10031\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44346\
        );

    \I__10030\ : Odrv4
    port map (
            O => \N__44352\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10029\ : Odrv4
    port map (
            O => \N__44349\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__44346\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__10027\ : CascadeMux
    port map (
            O => \N__44339\,
            I => \N__44336\
        );

    \I__10026\ : InMux
    port map (
            O => \N__44336\,
            I => \N__44329\
        );

    \I__10025\ : InMux
    port map (
            O => \N__44335\,
            I => \N__44329\
        );

    \I__10024\ : InMux
    port map (
            O => \N__44334\,
            I => \N__44326\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__44329\,
            I => \N__44323\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__44326\,
            I => \N__44318\
        );

    \I__10021\ : Span4Mux_v
    port map (
            O => \N__44323\,
            I => \N__44318\
        );

    \I__10020\ : Span4Mux_v
    port map (
            O => \N__44318\,
            I => \N__44314\
        );

    \I__10019\ : InMux
    port map (
            O => \N__44317\,
            I => \N__44311\
        );

    \I__10018\ : Odrv4
    port map (
            O => \N__44314\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__44311\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10016\ : CascadeMux
    port map (
            O => \N__44306\,
            I => \N__44303\
        );

    \I__10015\ : InMux
    port map (
            O => \N__44303\,
            I => \N__44300\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__44300\,
            I => \N__44297\
        );

    \I__10013\ : Odrv4
    port map (
            O => \N__44297\,
            I => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\
        );

    \I__10012\ : InMux
    port map (
            O => \N__44294\,
            I => \N__44291\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__44291\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__10010\ : CascadeMux
    port map (
            O => \N__44288\,
            I => \N__44285\
        );

    \I__10009\ : InMux
    port map (
            O => \N__44285\,
            I => \N__44282\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__44282\,
            I => \N__44279\
        );

    \I__10007\ : Odrv4
    port map (
            O => \N__44279\,
            I => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\
        );

    \I__10006\ : CascadeMux
    port map (
            O => \N__44276\,
            I => \N__44273\
        );

    \I__10005\ : InMux
    port map (
            O => \N__44273\,
            I => \N__44270\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__44270\,
            I => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\
        );

    \I__10003\ : CascadeMux
    port map (
            O => \N__44267\,
            I => \N__44264\
        );

    \I__10002\ : InMux
    port map (
            O => \N__44264\,
            I => \N__44259\
        );

    \I__10001\ : InMux
    port map (
            O => \N__44263\,
            I => \N__44256\
        );

    \I__10000\ : InMux
    port map (
            O => \N__44262\,
            I => \N__44253\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__44259\,
            I => \N__44250\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__44256\,
            I => \N__44247\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__44253\,
            I => \N__44244\
        );

    \I__9996\ : Span4Mux_h
    port map (
            O => \N__44250\,
            I => \N__44241\
        );

    \I__9995\ : Span4Mux_h
    port map (
            O => \N__44247\,
            I => \N__44238\
        );

    \I__9994\ : Span4Mux_h
    port map (
            O => \N__44244\,
            I => \N__44232\
        );

    \I__9993\ : Span4Mux_v
    port map (
            O => \N__44241\,
            I => \N__44232\
        );

    \I__9992\ : Span4Mux_v
    port map (
            O => \N__44238\,
            I => \N__44229\
        );

    \I__9991\ : InMux
    port map (
            O => \N__44237\,
            I => \N__44226\
        );

    \I__9990\ : Odrv4
    port map (
            O => \N__44232\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__9989\ : Odrv4
    port map (
            O => \N__44229\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__44226\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__9987\ : CascadeMux
    port map (
            O => \N__44219\,
            I => \N__44216\
        );

    \I__9986\ : InMux
    port map (
            O => \N__44216\,
            I => \N__44213\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__44213\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__9984\ : CascadeMux
    port map (
            O => \N__44210\,
            I => \N__44207\
        );

    \I__9983\ : InMux
    port map (
            O => \N__44207\,
            I => \N__44200\
        );

    \I__9982\ : InMux
    port map (
            O => \N__44206\,
            I => \N__44200\
        );

    \I__9981\ : InMux
    port map (
            O => \N__44205\,
            I => \N__44197\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__44200\,
            I => \N__44194\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__44197\,
            I => \N__44190\
        );

    \I__9978\ : Span12Mux_s10_h
    port map (
            O => \N__44194\,
            I => \N__44187\
        );

    \I__9977\ : InMux
    port map (
            O => \N__44193\,
            I => \N__44184\
        );

    \I__9976\ : Odrv4
    port map (
            O => \N__44190\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9975\ : Odrv12
    port map (
            O => \N__44187\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__44184\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9973\ : InMux
    port map (
            O => \N__44177\,
            I => \N__44174\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__44174\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__9971\ : CascadeMux
    port map (
            O => \N__44171\,
            I => \N__44168\
        );

    \I__9970\ : InMux
    port map (
            O => \N__44168\,
            I => \N__44162\
        );

    \I__9969\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44162\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__44162\,
            I => \N__44158\
        );

    \I__9967\ : InMux
    port map (
            O => \N__44161\,
            I => \N__44155\
        );

    \I__9966\ : Span4Mux_h
    port map (
            O => \N__44158\,
            I => \N__44152\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__44155\,
            I => \N__44146\
        );

    \I__9964\ : Span4Mux_v
    port map (
            O => \N__44152\,
            I => \N__44146\
        );

    \I__9963\ : InMux
    port map (
            O => \N__44151\,
            I => \N__44143\
        );

    \I__9962\ : Odrv4
    port map (
            O => \N__44146\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__44143\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9960\ : CascadeMux
    port map (
            O => \N__44138\,
            I => \N__44135\
        );

    \I__9959\ : InMux
    port map (
            O => \N__44135\,
            I => \N__44132\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__44132\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__9957\ : CascadeMux
    port map (
            O => \N__44129\,
            I => \N__44126\
        );

    \I__9956\ : InMux
    port map (
            O => \N__44126\,
            I => \N__44123\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__44123\,
            I => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\
        );

    \I__9954\ : InMux
    port map (
            O => \N__44120\,
            I => \N__44104\
        );

    \I__9953\ : InMux
    port map (
            O => \N__44119\,
            I => \N__44104\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44118\,
            I => \N__44104\
        );

    \I__9951\ : InMux
    port map (
            O => \N__44117\,
            I => \N__44104\
        );

    \I__9950\ : InMux
    port map (
            O => \N__44116\,
            I => \N__44095\
        );

    \I__9949\ : InMux
    port map (
            O => \N__44115\,
            I => \N__44095\
        );

    \I__9948\ : InMux
    port map (
            O => \N__44114\,
            I => \N__44095\
        );

    \I__9947\ : InMux
    port map (
            O => \N__44113\,
            I => \N__44095\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__44104\,
            I => \N__44072\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__44095\,
            I => \N__44072\
        );

    \I__9944\ : InMux
    port map (
            O => \N__44094\,
            I => \N__44063\
        );

    \I__9943\ : InMux
    port map (
            O => \N__44093\,
            I => \N__44063\
        );

    \I__9942\ : InMux
    port map (
            O => \N__44092\,
            I => \N__44063\
        );

    \I__9941\ : InMux
    port map (
            O => \N__44091\,
            I => \N__44063\
        );

    \I__9940\ : InMux
    port map (
            O => \N__44090\,
            I => \N__44058\
        );

    \I__9939\ : InMux
    port map (
            O => \N__44089\,
            I => \N__44058\
        );

    \I__9938\ : InMux
    port map (
            O => \N__44088\,
            I => \N__44045\
        );

    \I__9937\ : InMux
    port map (
            O => \N__44087\,
            I => \N__44045\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44045\
        );

    \I__9935\ : InMux
    port map (
            O => \N__44085\,
            I => \N__44045\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44084\,
            I => \N__44036\
        );

    \I__9933\ : InMux
    port map (
            O => \N__44083\,
            I => \N__44036\
        );

    \I__9932\ : InMux
    port map (
            O => \N__44082\,
            I => \N__44036\
        );

    \I__9931\ : InMux
    port map (
            O => \N__44081\,
            I => \N__44036\
        );

    \I__9930\ : InMux
    port map (
            O => \N__44080\,
            I => \N__44027\
        );

    \I__9929\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44027\
        );

    \I__9928\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44027\
        );

    \I__9927\ : InMux
    port map (
            O => \N__44077\,
            I => \N__44027\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__44072\,
            I => \N__44020\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__44063\,
            I => \N__44020\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__44058\,
            I => \N__44020\
        );

    \I__9923\ : InMux
    port map (
            O => \N__44057\,
            I => \N__44011\
        );

    \I__9922\ : InMux
    port map (
            O => \N__44056\,
            I => \N__44011\
        );

    \I__9921\ : InMux
    port map (
            O => \N__44055\,
            I => \N__44011\
        );

    \I__9920\ : InMux
    port map (
            O => \N__44054\,
            I => \N__44011\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__44045\,
            I => \N__44006\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__44036\,
            I => \N__44006\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__44027\,
            I => \N__44001\
        );

    \I__9916\ : Span4Mux_v
    port map (
            O => \N__44020\,
            I => \N__44001\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__44011\,
            I => \N__43998\
        );

    \I__9914\ : Span4Mux_v
    port map (
            O => \N__44006\,
            I => \N__43993\
        );

    \I__9913\ : Span4Mux_h
    port map (
            O => \N__44001\,
            I => \N__43993\
        );

    \I__9912\ : Odrv4
    port map (
            O => \N__43998\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9911\ : Odrv4
    port map (
            O => \N__43993\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9910\ : InMux
    port map (
            O => \N__43988\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__9909\ : InMux
    port map (
            O => \N__43985\,
            I => \N__43981\
        );

    \I__9908\ : InMux
    port map (
            O => \N__43984\,
            I => \N__43978\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__43981\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__43978\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__9905\ : CEMux
    port map (
            O => \N__43973\,
            I => \N__43970\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__43970\,
            I => \N__43966\
        );

    \I__9903\ : CEMux
    port map (
            O => \N__43969\,
            I => \N__43962\
        );

    \I__9902\ : Span4Mux_v
    port map (
            O => \N__43966\,
            I => \N__43959\
        );

    \I__9901\ : CEMux
    port map (
            O => \N__43965\,
            I => \N__43956\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__43962\,
            I => \N__43948\
        );

    \I__9899\ : Span4Mux_h
    port map (
            O => \N__43959\,
            I => \N__43948\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__43956\,
            I => \N__43948\
        );

    \I__9897\ : CEMux
    port map (
            O => \N__43955\,
            I => \N__43945\
        );

    \I__9896\ : Sp12to4
    port map (
            O => \N__43948\,
            I => \N__43940\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__43945\,
            I => \N__43940\
        );

    \I__9894\ : Odrv12
    port map (
            O => \N__43940\,
            I => \delay_measurement_inst.delay_tr_timer.N_305_i\
        );

    \I__9893\ : InMux
    port map (
            O => \N__43937\,
            I => \N__43934\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__43934\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__9891\ : InMux
    port map (
            O => \N__43931\,
            I => \N__43927\
        );

    \I__9890\ : InMux
    port map (
            O => \N__43930\,
            I => \N__43924\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__43927\,
            I => \N__43921\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__43924\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9887\ : Odrv12
    port map (
            O => \N__43921\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9886\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43911\
        );

    \I__9885\ : InMux
    port map (
            O => \N__43915\,
            I => \N__43908\
        );

    \I__9884\ : InMux
    port map (
            O => \N__43914\,
            I => \N__43905\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__43911\,
            I => \N__43900\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__43908\,
            I => \N__43900\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__43905\,
            I => \N__43895\
        );

    \I__9880\ : Span4Mux_v
    port map (
            O => \N__43900\,
            I => \N__43895\
        );

    \I__9879\ : Odrv4
    port map (
            O => \N__43895\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__9878\ : CascadeMux
    port map (
            O => \N__43892\,
            I => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\
        );

    \I__9877\ : InMux
    port map (
            O => \N__43889\,
            I => \N__43886\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__43886\,
            I => \N__43883\
        );

    \I__9875\ : Span4Mux_h
    port map (
            O => \N__43883\,
            I => \N__43875\
        );

    \I__9874\ : InMux
    port map (
            O => \N__43882\,
            I => \N__43872\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43863\
        );

    \I__9872\ : InMux
    port map (
            O => \N__43880\,
            I => \N__43863\
        );

    \I__9871\ : InMux
    port map (
            O => \N__43879\,
            I => \N__43863\
        );

    \I__9870\ : InMux
    port map (
            O => \N__43878\,
            I => \N__43863\
        );

    \I__9869\ : Odrv4
    port map (
            O => \N__43875\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__43872\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__43863\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9866\ : InMux
    port map (
            O => \N__43856\,
            I => \N__43852\
        );

    \I__9865\ : InMux
    port map (
            O => \N__43855\,
            I => \N__43849\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__43852\,
            I => \N__43846\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__43849\,
            I => \N__43843\
        );

    \I__9862\ : Span4Mux_h
    port map (
            O => \N__43846\,
            I => \N__43840\
        );

    \I__9861\ : Span4Mux_h
    port map (
            O => \N__43843\,
            I => \N__43837\
        );

    \I__9860\ : Span4Mux_v
    port map (
            O => \N__43840\,
            I => \N__43834\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__43837\,
            I => \N__43831\
        );

    \I__9858\ : Odrv4
    port map (
            O => \N__43834\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__9857\ : Odrv4
    port map (
            O => \N__43831\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__9856\ : InMux
    port map (
            O => \N__43826\,
            I => \N__43808\
        );

    \I__9855\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43808\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43824\,
            I => \N__43808\
        );

    \I__9853\ : CascadeMux
    port map (
            O => \N__43823\,
            I => \N__43805\
        );

    \I__9852\ : CascadeMux
    port map (
            O => \N__43822\,
            I => \N__43801\
        );

    \I__9851\ : InMux
    port map (
            O => \N__43821\,
            I => \N__43779\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43779\
        );

    \I__9849\ : InMux
    port map (
            O => \N__43819\,
            I => \N__43779\
        );

    \I__9848\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43779\
        );

    \I__9847\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43779\
        );

    \I__9846\ : InMux
    port map (
            O => \N__43816\,
            I => \N__43779\
        );

    \I__9845\ : InMux
    port map (
            O => \N__43815\,
            I => \N__43779\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__43808\,
            I => \N__43772\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43805\,
            I => \N__43767\
        );

    \I__9842\ : InMux
    port map (
            O => \N__43804\,
            I => \N__43767\
        );

    \I__9841\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43750\
        );

    \I__9840\ : InMux
    port map (
            O => \N__43800\,
            I => \N__43750\
        );

    \I__9839\ : InMux
    port map (
            O => \N__43799\,
            I => \N__43750\
        );

    \I__9838\ : InMux
    port map (
            O => \N__43798\,
            I => \N__43750\
        );

    \I__9837\ : InMux
    port map (
            O => \N__43797\,
            I => \N__43750\
        );

    \I__9836\ : InMux
    port map (
            O => \N__43796\,
            I => \N__43750\
        );

    \I__9835\ : InMux
    port map (
            O => \N__43795\,
            I => \N__43750\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43794\,
            I => \N__43750\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__43779\,
            I => \N__43747\
        );

    \I__9832\ : InMux
    port map (
            O => \N__43778\,
            I => \N__43738\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43777\,
            I => \N__43738\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43776\,
            I => \N__43738\
        );

    \I__9829\ : InMux
    port map (
            O => \N__43775\,
            I => \N__43738\
        );

    \I__9828\ : Span4Mux_v
    port map (
            O => \N__43772\,
            I => \N__43735\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__43767\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9826\ : LocalMux
    port map (
            O => \N__43750\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9825\ : Odrv4
    port map (
            O => \N__43747\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__43738\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9823\ : Odrv4
    port map (
            O => \N__43735\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__9822\ : CascadeMux
    port map (
            O => \N__43724\,
            I => \N__43713\
        );

    \I__9821\ : CascadeMux
    port map (
            O => \N__43723\,
            I => \N__43709\
        );

    \I__9820\ : CascadeMux
    port map (
            O => \N__43722\,
            I => \N__43705\
        );

    \I__9819\ : CascadeMux
    port map (
            O => \N__43721\,
            I => \N__43701\
        );

    \I__9818\ : CascadeMux
    port map (
            O => \N__43720\,
            I => \N__43697\
        );

    \I__9817\ : CascadeMux
    port map (
            O => \N__43719\,
            I => \N__43692\
        );

    \I__9816\ : CascadeMux
    port map (
            O => \N__43718\,
            I => \N__43688\
        );

    \I__9815\ : CascadeMux
    port map (
            O => \N__43717\,
            I => \N__43684\
        );

    \I__9814\ : InMux
    port map (
            O => \N__43716\,
            I => \N__43678\
        );

    \I__9813\ : InMux
    port map (
            O => \N__43713\,
            I => \N__43678\
        );

    \I__9812\ : InMux
    port map (
            O => \N__43712\,
            I => \N__43661\
        );

    \I__9811\ : InMux
    port map (
            O => \N__43709\,
            I => \N__43661\
        );

    \I__9810\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43661\
        );

    \I__9809\ : InMux
    port map (
            O => \N__43705\,
            I => \N__43661\
        );

    \I__9808\ : InMux
    port map (
            O => \N__43704\,
            I => \N__43661\
        );

    \I__9807\ : InMux
    port map (
            O => \N__43701\,
            I => \N__43661\
        );

    \I__9806\ : InMux
    port map (
            O => \N__43700\,
            I => \N__43661\
        );

    \I__9805\ : InMux
    port map (
            O => \N__43697\,
            I => \N__43661\
        );

    \I__9804\ : InMux
    port map (
            O => \N__43696\,
            I => \N__43657\
        );

    \I__9803\ : InMux
    port map (
            O => \N__43695\,
            I => \N__43644\
        );

    \I__9802\ : InMux
    port map (
            O => \N__43692\,
            I => \N__43644\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43691\,
            I => \N__43644\
        );

    \I__9800\ : InMux
    port map (
            O => \N__43688\,
            I => \N__43644\
        );

    \I__9799\ : InMux
    port map (
            O => \N__43687\,
            I => \N__43644\
        );

    \I__9798\ : InMux
    port map (
            O => \N__43684\,
            I => \N__43644\
        );

    \I__9797\ : CascadeMux
    port map (
            O => \N__43683\,
            I => \N__43641\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__43678\,
            I => \N__43635\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__43661\,
            I => \N__43635\
        );

    \I__9794\ : CascadeMux
    port map (
            O => \N__43660\,
            I => \N__43631\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__43657\,
            I => \N__43624\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__43644\,
            I => \N__43624\
        );

    \I__9791\ : InMux
    port map (
            O => \N__43641\,
            I => \N__43619\
        );

    \I__9790\ : InMux
    port map (
            O => \N__43640\,
            I => \N__43619\
        );

    \I__9789\ : Span4Mux_v
    port map (
            O => \N__43635\,
            I => \N__43616\
        );

    \I__9788\ : InMux
    port map (
            O => \N__43634\,
            I => \N__43607\
        );

    \I__9787\ : InMux
    port map (
            O => \N__43631\,
            I => \N__43607\
        );

    \I__9786\ : InMux
    port map (
            O => \N__43630\,
            I => \N__43607\
        );

    \I__9785\ : InMux
    port map (
            O => \N__43629\,
            I => \N__43607\
        );

    \I__9784\ : Span4Mux_h
    port map (
            O => \N__43624\,
            I => \N__43602\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43619\,
            I => \N__43602\
        );

    \I__9782\ : Sp12to4
    port map (
            O => \N__43616\,
            I => \N__43596\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__43607\,
            I => \N__43596\
        );

    \I__9780\ : Span4Mux_v
    port map (
            O => \N__43602\,
            I => \N__43593\
        );

    \I__9779\ : InMux
    port map (
            O => \N__43601\,
            I => \N__43590\
        );

    \I__9778\ : Span12Mux_h
    port map (
            O => \N__43596\,
            I => \N__43587\
        );

    \I__9777\ : Span4Mux_h
    port map (
            O => \N__43593\,
            I => \N__43584\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__43590\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9775\ : Odrv12
    port map (
            O => \N__43587\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9774\ : Odrv4
    port map (
            O => \N__43584\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__9773\ : CascadeMux
    port map (
            O => \N__43577\,
            I => \N__43572\
        );

    \I__9772\ : CascadeMux
    port map (
            O => \N__43576\,
            I => \N__43569\
        );

    \I__9771\ : CascadeMux
    port map (
            O => \N__43575\,
            I => \N__43566\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43572\,
            I => \N__43547\
        );

    \I__9769\ : InMux
    port map (
            O => \N__43569\,
            I => \N__43547\
        );

    \I__9768\ : InMux
    port map (
            O => \N__43566\,
            I => \N__43547\
        );

    \I__9767\ : InMux
    port map (
            O => \N__43565\,
            I => \N__43538\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43564\,
            I => \N__43538\
        );

    \I__9765\ : InMux
    port map (
            O => \N__43563\,
            I => \N__43538\
        );

    \I__9764\ : InMux
    port map (
            O => \N__43562\,
            I => \N__43538\
        );

    \I__9763\ : InMux
    port map (
            O => \N__43561\,
            I => \N__43533\
        );

    \I__9762\ : InMux
    port map (
            O => \N__43560\,
            I => \N__43533\
        );

    \I__9761\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43530\
        );

    \I__9760\ : CascadeMux
    port map (
            O => \N__43558\,
            I => \N__43527\
        );

    \I__9759\ : CascadeMux
    port map (
            O => \N__43557\,
            I => \N__43523\
        );

    \I__9758\ : CascadeMux
    port map (
            O => \N__43556\,
            I => \N__43520\
        );

    \I__9757\ : CascadeMux
    port map (
            O => \N__43555\,
            I => \N__43510\
        );

    \I__9756\ : CascadeMux
    port map (
            O => \N__43554\,
            I => \N__43507\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__43547\,
            I => \N__43497\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__43538\,
            I => \N__43497\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__43533\,
            I => \N__43497\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__43530\,
            I => \N__43497\
        );

    \I__9751\ : InMux
    port map (
            O => \N__43527\,
            I => \N__43488\
        );

    \I__9750\ : InMux
    port map (
            O => \N__43526\,
            I => \N__43488\
        );

    \I__9749\ : InMux
    port map (
            O => \N__43523\,
            I => \N__43488\
        );

    \I__9748\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43488\
        );

    \I__9747\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43483\
        );

    \I__9746\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43483\
        );

    \I__9745\ : InMux
    port map (
            O => \N__43517\,
            I => \N__43480\
        );

    \I__9744\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43471\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43515\,
            I => \N__43471\
        );

    \I__9742\ : InMux
    port map (
            O => \N__43514\,
            I => \N__43471\
        );

    \I__9741\ : InMux
    port map (
            O => \N__43513\,
            I => \N__43471\
        );

    \I__9740\ : InMux
    port map (
            O => \N__43510\,
            I => \N__43464\
        );

    \I__9739\ : InMux
    port map (
            O => \N__43507\,
            I => \N__43464\
        );

    \I__9738\ : InMux
    port map (
            O => \N__43506\,
            I => \N__43464\
        );

    \I__9737\ : Span4Mux_h
    port map (
            O => \N__43497\,
            I => \N__43461\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__43488\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__43483\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__43480\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__43471\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__43464\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__9731\ : Odrv4
    port map (
            O => \N__43461\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__9730\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43445\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__43445\,
            I => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__9728\ : InMux
    port map (
            O => \N__43442\,
            I => \N__43439\
        );

    \I__9727\ : LocalMux
    port map (
            O => \N__43439\,
            I => \N__43436\
        );

    \I__9726\ : Span4Mux_v
    port map (
            O => \N__43436\,
            I => \N__43432\
        );

    \I__9725\ : InMux
    port map (
            O => \N__43435\,
            I => \N__43429\
        );

    \I__9724\ : Span4Mux_v
    port map (
            O => \N__43432\,
            I => \N__43426\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__43429\,
            I => \N__43423\
        );

    \I__9722\ : Span4Mux_v
    port map (
            O => \N__43426\,
            I => \N__43420\
        );

    \I__9721\ : Span12Mux_h
    port map (
            O => \N__43423\,
            I => \N__43416\
        );

    \I__9720\ : Span4Mux_v
    port map (
            O => \N__43420\,
            I => \N__43413\
        );

    \I__9719\ : InMux
    port map (
            O => \N__43419\,
            I => \N__43410\
        );

    \I__9718\ : Odrv12
    port map (
            O => \N__43416\,
            I => \il_min_comp1_D2\
        );

    \I__9717\ : Odrv4
    port map (
            O => \N__43413\,
            I => \il_min_comp1_D2\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__43410\,
            I => \il_min_comp1_D2\
        );

    \I__9715\ : InMux
    port map (
            O => \N__43403\,
            I => \N__43398\
        );

    \I__9714\ : InMux
    port map (
            O => \N__43402\,
            I => \N__43393\
        );

    \I__9713\ : InMux
    port map (
            O => \N__43401\,
            I => \N__43393\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__43398\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__43393\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__9710\ : CascadeMux
    port map (
            O => \N__43388\,
            I => \N__43385\
        );

    \I__9709\ : InMux
    port map (
            O => \N__43385\,
            I => \N__43382\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__43382\,
            I => \N__43377\
        );

    \I__9707\ : InMux
    port map (
            O => \N__43381\,
            I => \N__43374\
        );

    \I__9706\ : InMux
    port map (
            O => \N__43380\,
            I => \N__43371\
        );

    \I__9705\ : Span4Mux_v
    port map (
            O => \N__43377\,
            I => \N__43368\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__43374\,
            I => \N__43364\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__43371\,
            I => \N__43361\
        );

    \I__9702\ : Span4Mux_v
    port map (
            O => \N__43368\,
            I => \N__43358\
        );

    \I__9701\ : CascadeMux
    port map (
            O => \N__43367\,
            I => \N__43355\
        );

    \I__9700\ : Span12Mux_s7_v
    port map (
            O => \N__43364\,
            I => \N__43352\
        );

    \I__9699\ : Span4Mux_v
    port map (
            O => \N__43361\,
            I => \N__43347\
        );

    \I__9698\ : Span4Mux_h
    port map (
            O => \N__43358\,
            I => \N__43347\
        );

    \I__9697\ : InMux
    port map (
            O => \N__43355\,
            I => \N__43344\
        );

    \I__9696\ : Span12Mux_v
    port map (
            O => \N__43352\,
            I => \N__43341\
        );

    \I__9695\ : Odrv4
    port map (
            O => \N__43347\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9694\ : LocalMux
    port map (
            O => \N__43344\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9693\ : Odrv12
    port map (
            O => \N__43341\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9692\ : InMux
    port map (
            O => \N__43334\,
            I => \N__43330\
        );

    \I__9691\ : InMux
    port map (
            O => \N__43333\,
            I => \N__43327\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__43330\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__43327\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__9688\ : InMux
    port map (
            O => \N__43322\,
            I => \N__43317\
        );

    \I__9687\ : InMux
    port map (
            O => \N__43321\,
            I => \N__43312\
        );

    \I__9686\ : InMux
    port map (
            O => \N__43320\,
            I => \N__43312\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__43317\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__43312\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__9683\ : InMux
    port map (
            O => \N__43307\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__9682\ : InMux
    port map (
            O => \N__43304\,
            I => \N__43299\
        );

    \I__9681\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43294\
        );

    \I__9680\ : InMux
    port map (
            O => \N__43302\,
            I => \N__43294\
        );

    \I__9679\ : LocalMux
    port map (
            O => \N__43299\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__43294\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__9677\ : InMux
    port map (
            O => \N__43289\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__9676\ : CascadeMux
    port map (
            O => \N__43286\,
            I => \N__43281\
        );

    \I__9675\ : CascadeMux
    port map (
            O => \N__43285\,
            I => \N__43278\
        );

    \I__9674\ : InMux
    port map (
            O => \N__43284\,
            I => \N__43275\
        );

    \I__9673\ : InMux
    port map (
            O => \N__43281\,
            I => \N__43270\
        );

    \I__9672\ : InMux
    port map (
            O => \N__43278\,
            I => \N__43270\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__43275\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__43270\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__9669\ : InMux
    port map (
            O => \N__43265\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__9668\ : CascadeMux
    port map (
            O => \N__43262\,
            I => \N__43257\
        );

    \I__9667\ : CascadeMux
    port map (
            O => \N__43261\,
            I => \N__43254\
        );

    \I__9666\ : InMux
    port map (
            O => \N__43260\,
            I => \N__43251\
        );

    \I__9665\ : InMux
    port map (
            O => \N__43257\,
            I => \N__43246\
        );

    \I__9664\ : InMux
    port map (
            O => \N__43254\,
            I => \N__43246\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__43251\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9662\ : LocalMux
    port map (
            O => \N__43246\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9661\ : InMux
    port map (
            O => \N__43241\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__9660\ : InMux
    port map (
            O => \N__43238\,
            I => \N__43233\
        );

    \I__9659\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43230\
        );

    \I__9658\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43227\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__43233\,
            I => \N__43224\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__43230\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__43227\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__9654\ : Odrv4
    port map (
            O => \N__43224\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__9653\ : InMux
    port map (
            O => \N__43217\,
            I => \bfn_17_10_0_\
        );

    \I__9652\ : InMux
    port map (
            O => \N__43214\,
            I => \N__43209\
        );

    \I__9651\ : InMux
    port map (
            O => \N__43213\,
            I => \N__43206\
        );

    \I__9650\ : InMux
    port map (
            O => \N__43212\,
            I => \N__43203\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__43209\,
            I => \N__43200\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__43206\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__43203\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9646\ : Odrv4
    port map (
            O => \N__43200\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__9645\ : InMux
    port map (
            O => \N__43193\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__9644\ : CascadeMux
    port map (
            O => \N__43190\,
            I => \N__43185\
        );

    \I__9643\ : CascadeMux
    port map (
            O => \N__43189\,
            I => \N__43182\
        );

    \I__9642\ : InMux
    port map (
            O => \N__43188\,
            I => \N__43179\
        );

    \I__9641\ : InMux
    port map (
            O => \N__43185\,
            I => \N__43174\
        );

    \I__9640\ : InMux
    port map (
            O => \N__43182\,
            I => \N__43174\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__43179\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__43174\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__9637\ : InMux
    port map (
            O => \N__43169\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__9636\ : CascadeMux
    port map (
            O => \N__43166\,
            I => \N__43161\
        );

    \I__9635\ : CascadeMux
    port map (
            O => \N__43165\,
            I => \N__43158\
        );

    \I__9634\ : InMux
    port map (
            O => \N__43164\,
            I => \N__43155\
        );

    \I__9633\ : InMux
    port map (
            O => \N__43161\,
            I => \N__43150\
        );

    \I__9632\ : InMux
    port map (
            O => \N__43158\,
            I => \N__43150\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__43155\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__43150\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__9629\ : InMux
    port map (
            O => \N__43145\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__9628\ : InMux
    port map (
            O => \N__43142\,
            I => \N__43138\
        );

    \I__9627\ : InMux
    port map (
            O => \N__43141\,
            I => \N__43135\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__43138\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__43135\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__9624\ : InMux
    port map (
            O => \N__43130\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__9623\ : InMux
    port map (
            O => \N__43127\,
            I => \N__43122\
        );

    \I__9622\ : InMux
    port map (
            O => \N__43126\,
            I => \N__43117\
        );

    \I__9621\ : InMux
    port map (
            O => \N__43125\,
            I => \N__43117\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__43122\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__43117\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__9618\ : InMux
    port map (
            O => \N__43112\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__9617\ : InMux
    port map (
            O => \N__43109\,
            I => \N__43104\
        );

    \I__9616\ : InMux
    port map (
            O => \N__43108\,
            I => \N__43099\
        );

    \I__9615\ : InMux
    port map (
            O => \N__43107\,
            I => \N__43099\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__43104\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__43099\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__9612\ : InMux
    port map (
            O => \N__43094\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__9611\ : CascadeMux
    port map (
            O => \N__43091\,
            I => \N__43086\
        );

    \I__9610\ : CascadeMux
    port map (
            O => \N__43090\,
            I => \N__43083\
        );

    \I__9609\ : InMux
    port map (
            O => \N__43089\,
            I => \N__43080\
        );

    \I__9608\ : InMux
    port map (
            O => \N__43086\,
            I => \N__43075\
        );

    \I__9607\ : InMux
    port map (
            O => \N__43083\,
            I => \N__43075\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__43080\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__43075\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__9604\ : InMux
    port map (
            O => \N__43070\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__9603\ : CascadeMux
    port map (
            O => \N__43067\,
            I => \N__43062\
        );

    \I__9602\ : CascadeMux
    port map (
            O => \N__43066\,
            I => \N__43059\
        );

    \I__9601\ : InMux
    port map (
            O => \N__43065\,
            I => \N__43056\
        );

    \I__9600\ : InMux
    port map (
            O => \N__43062\,
            I => \N__43051\
        );

    \I__9599\ : InMux
    port map (
            O => \N__43059\,
            I => \N__43051\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__43056\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__43051\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__9596\ : InMux
    port map (
            O => \N__43046\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__9595\ : InMux
    port map (
            O => \N__43043\,
            I => \N__43038\
        );

    \I__9594\ : InMux
    port map (
            O => \N__43042\,
            I => \N__43035\
        );

    \I__9593\ : InMux
    port map (
            O => \N__43041\,
            I => \N__43032\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__43038\,
            I => \N__43029\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__43035\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__43032\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__43029\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__9588\ : InMux
    port map (
            O => \N__43022\,
            I => \bfn_17_9_0_\
        );

    \I__9587\ : InMux
    port map (
            O => \N__43019\,
            I => \N__43014\
        );

    \I__9586\ : InMux
    port map (
            O => \N__43018\,
            I => \N__43011\
        );

    \I__9585\ : InMux
    port map (
            O => \N__43017\,
            I => \N__43008\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__43014\,
            I => \N__43005\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__43011\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__43008\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9581\ : Odrv4
    port map (
            O => \N__43005\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9580\ : InMux
    port map (
            O => \N__42998\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__9579\ : CascadeMux
    port map (
            O => \N__42995\,
            I => \N__42990\
        );

    \I__9578\ : CascadeMux
    port map (
            O => \N__42994\,
            I => \N__42987\
        );

    \I__9577\ : InMux
    port map (
            O => \N__42993\,
            I => \N__42984\
        );

    \I__9576\ : InMux
    port map (
            O => \N__42990\,
            I => \N__42979\
        );

    \I__9575\ : InMux
    port map (
            O => \N__42987\,
            I => \N__42979\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__42984\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__42979\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__9572\ : InMux
    port map (
            O => \N__42974\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__9571\ : CascadeMux
    port map (
            O => \N__42971\,
            I => \N__42966\
        );

    \I__9570\ : CascadeMux
    port map (
            O => \N__42970\,
            I => \N__42963\
        );

    \I__9569\ : InMux
    port map (
            O => \N__42969\,
            I => \N__42960\
        );

    \I__9568\ : InMux
    port map (
            O => \N__42966\,
            I => \N__42955\
        );

    \I__9567\ : InMux
    port map (
            O => \N__42963\,
            I => \N__42955\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__42960\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__42955\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__9564\ : InMux
    port map (
            O => \N__42950\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__9563\ : InMux
    port map (
            O => \N__42947\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__9562\ : InMux
    port map (
            O => \N__42944\,
            I => \N__42939\
        );

    \I__9561\ : InMux
    port map (
            O => \N__42943\,
            I => \N__42934\
        );

    \I__9560\ : InMux
    port map (
            O => \N__42942\,
            I => \N__42934\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__42939\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__42934\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__9557\ : InMux
    port map (
            O => \N__42929\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__9556\ : InMux
    port map (
            O => \N__42926\,
            I => \N__42921\
        );

    \I__9555\ : InMux
    port map (
            O => \N__42925\,
            I => \N__42916\
        );

    \I__9554\ : InMux
    port map (
            O => \N__42924\,
            I => \N__42916\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__42921\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__42916\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__9551\ : InMux
    port map (
            O => \N__42911\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__9550\ : CascadeMux
    port map (
            O => \N__42908\,
            I => \N__42903\
        );

    \I__9549\ : CascadeMux
    port map (
            O => \N__42907\,
            I => \N__42900\
        );

    \I__9548\ : InMux
    port map (
            O => \N__42906\,
            I => \N__42897\
        );

    \I__9547\ : InMux
    port map (
            O => \N__42903\,
            I => \N__42892\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42900\,
            I => \N__42892\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__42897\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__42892\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__9543\ : InMux
    port map (
            O => \N__42887\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__9542\ : CascadeMux
    port map (
            O => \N__42884\,
            I => \N__42879\
        );

    \I__9541\ : CascadeMux
    port map (
            O => \N__42883\,
            I => \N__42876\
        );

    \I__9540\ : InMux
    port map (
            O => \N__42882\,
            I => \N__42873\
        );

    \I__9539\ : InMux
    port map (
            O => \N__42879\,
            I => \N__42868\
        );

    \I__9538\ : InMux
    port map (
            O => \N__42876\,
            I => \N__42868\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__42873\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__42868\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42863\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__9534\ : InMux
    port map (
            O => \N__42860\,
            I => \N__42855\
        );

    \I__9533\ : InMux
    port map (
            O => \N__42859\,
            I => \N__42852\
        );

    \I__9532\ : InMux
    port map (
            O => \N__42858\,
            I => \N__42849\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__42855\,
            I => \N__42846\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__42852\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__42849\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__9528\ : Odrv4
    port map (
            O => \N__42846\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__9527\ : InMux
    port map (
            O => \N__42839\,
            I => \bfn_17_8_0_\
        );

    \I__9526\ : InMux
    port map (
            O => \N__42836\,
            I => \N__42831\
        );

    \I__9525\ : InMux
    port map (
            O => \N__42835\,
            I => \N__42828\
        );

    \I__9524\ : InMux
    port map (
            O => \N__42834\,
            I => \N__42825\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__42831\,
            I => \N__42822\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__42828\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__42825\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__9520\ : Odrv4
    port map (
            O => \N__42822\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__9519\ : InMux
    port map (
            O => \N__42815\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__9518\ : CascadeMux
    port map (
            O => \N__42812\,
            I => \N__42807\
        );

    \I__9517\ : CascadeMux
    port map (
            O => \N__42811\,
            I => \N__42804\
        );

    \I__9516\ : InMux
    port map (
            O => \N__42810\,
            I => \N__42801\
        );

    \I__9515\ : InMux
    port map (
            O => \N__42807\,
            I => \N__42796\
        );

    \I__9514\ : InMux
    port map (
            O => \N__42804\,
            I => \N__42796\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__42801\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__42796\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42791\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__9510\ : CascadeMux
    port map (
            O => \N__42788\,
            I => \N__42783\
        );

    \I__9509\ : CascadeMux
    port map (
            O => \N__42787\,
            I => \N__42780\
        );

    \I__9508\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42777\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42783\,
            I => \N__42772\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42780\,
            I => \N__42772\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__42777\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__42772\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42767\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42764\,
            I => \N__42761\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42761\,
            I => \N__42757\
        );

    \I__9500\ : InMux
    port map (
            O => \N__42760\,
            I => \N__42754\
        );

    \I__9499\ : Span4Mux_v
    port map (
            O => \N__42757\,
            I => \N__42751\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42754\,
            I => \N__42748\
        );

    \I__9497\ : Span4Mux_v
    port map (
            O => \N__42751\,
            I => \N__42741\
        );

    \I__9496\ : Span4Mux_h
    port map (
            O => \N__42748\,
            I => \N__42741\
        );

    \I__9495\ : InMux
    port map (
            O => \N__42747\,
            I => \N__42738\
        );

    \I__9494\ : InMux
    port map (
            O => \N__42746\,
            I => \N__42735\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__42741\,
            I => measured_delay_tr_16
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__42738\,
            I => measured_delay_tr_16
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__42735\,
            I => measured_delay_tr_16
        );

    \I__9490\ : CascadeMux
    port map (
            O => \N__42728\,
            I => \N__42725\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42725\,
            I => \N__42722\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__42722\,
            I => \N__42719\
        );

    \I__9487\ : Span4Mux_v
    port map (
            O => \N__42719\,
            I => \N__42716\
        );

    \I__9486\ : Span4Mux_h
    port map (
            O => \N__42716\,
            I => \N__42713\
        );

    \I__9485\ : Odrv4
    port map (
            O => \N__42713\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__9484\ : CEMux
    port map (
            O => \N__42710\,
            I => \N__42706\
        );

    \I__9483\ : CEMux
    port map (
            O => \N__42709\,
            I => \N__42702\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__42706\,
            I => \N__42697\
        );

    \I__9481\ : CEMux
    port map (
            O => \N__42705\,
            I => \N__42694\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__42702\,
            I => \N__42691\
        );

    \I__9479\ : CEMux
    port map (
            O => \N__42701\,
            I => \N__42688\
        );

    \I__9478\ : CEMux
    port map (
            O => \N__42700\,
            I => \N__42684\
        );

    \I__9477\ : Span4Mux_v
    port map (
            O => \N__42697\,
            I => \N__42680\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__42694\,
            I => \N__42673\
        );

    \I__9475\ : Span4Mux_v
    port map (
            O => \N__42691\,
            I => \N__42673\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__42688\,
            I => \N__42673\
        );

    \I__9473\ : CEMux
    port map (
            O => \N__42687\,
            I => \N__42670\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__42684\,
            I => \N__42667\
        );

    \I__9471\ : CEMux
    port map (
            O => \N__42683\,
            I => \N__42664\
        );

    \I__9470\ : Span4Mux_h
    port map (
            O => \N__42680\,
            I => \N__42659\
        );

    \I__9469\ : Span4Mux_v
    port map (
            O => \N__42673\,
            I => \N__42659\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__42670\,
            I => \N__42656\
        );

    \I__9467\ : Span4Mux_h
    port map (
            O => \N__42667\,
            I => \N__42653\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__42664\,
            I => \N__42650\
        );

    \I__9465\ : Odrv4
    port map (
            O => \N__42659\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9464\ : Odrv12
    port map (
            O => \N__42656\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9463\ : Odrv4
    port map (
            O => \N__42653\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9462\ : Odrv12
    port map (
            O => \N__42650\,
            I => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9461\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42638\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__42638\,
            I => \N__42635\
        );

    \I__9459\ : Span4Mux_h
    port map (
            O => \N__42635\,
            I => \N__42631\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42634\,
            I => \N__42628\
        );

    \I__9457\ : Span4Mux_h
    port map (
            O => \N__42631\,
            I => \N__42625\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__42628\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__9455\ : Odrv4
    port map (
            O => \N__42625\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__9454\ : InMux
    port map (
            O => \N__42620\,
            I => \N__42617\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__42617\,
            I => \N__42613\
        );

    \I__9452\ : InMux
    port map (
            O => \N__42616\,
            I => \N__42610\
        );

    \I__9451\ : Span4Mux_h
    port map (
            O => \N__42613\,
            I => \N__42607\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__42610\,
            I => \N__42603\
        );

    \I__9449\ : Span4Mux_v
    port map (
            O => \N__42607\,
            I => \N__42600\
        );

    \I__9448\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42597\
        );

    \I__9447\ : Odrv4
    port map (
            O => \N__42603\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__9446\ : Odrv4
    port map (
            O => \N__42600\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__42597\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__9444\ : InMux
    port map (
            O => \N__42590\,
            I => \N__42586\
        );

    \I__9443\ : InMux
    port map (
            O => \N__42589\,
            I => \N__42583\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__42586\,
            I => \N__42578\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__42583\,
            I => \N__42575\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42582\,
            I => \N__42572\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42581\,
            I => \N__42569\
        );

    \I__9438\ : Span12Mux_h
    port map (
            O => \N__42578\,
            I => \N__42566\
        );

    \I__9437\ : Span4Mux_v
    port map (
            O => \N__42575\,
            I => \N__42563\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__42572\,
            I => \N__42560\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__42569\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__9434\ : Odrv12
    port map (
            O => \N__42566\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__9433\ : Odrv4
    port map (
            O => \N__42563\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__42560\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__9431\ : InMux
    port map (
            O => \N__42551\,
            I => \bfn_17_7_0_\
        );

    \I__9430\ : InMux
    port map (
            O => \N__42548\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__9429\ : CascadeMux
    port map (
            O => \N__42545\,
            I => \N__42540\
        );

    \I__9428\ : CascadeMux
    port map (
            O => \N__42544\,
            I => \N__42537\
        );

    \I__9427\ : InMux
    port map (
            O => \N__42543\,
            I => \N__42534\
        );

    \I__9426\ : InMux
    port map (
            O => \N__42540\,
            I => \N__42529\
        );

    \I__9425\ : InMux
    port map (
            O => \N__42537\,
            I => \N__42529\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__42534\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__42529\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42524\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__9421\ : CascadeMux
    port map (
            O => \N__42521\,
            I => \N__42516\
        );

    \I__9420\ : CascadeMux
    port map (
            O => \N__42520\,
            I => \N__42513\
        );

    \I__9419\ : InMux
    port map (
            O => \N__42519\,
            I => \N__42510\
        );

    \I__9418\ : InMux
    port map (
            O => \N__42516\,
            I => \N__42505\
        );

    \I__9417\ : InMux
    port map (
            O => \N__42513\,
            I => \N__42505\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__42510\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__42505\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__9414\ : CascadeMux
    port map (
            O => \N__42500\,
            I => \N__42496\
        );

    \I__9413\ : CascadeMux
    port map (
            O => \N__42499\,
            I => \N__42493\
        );

    \I__9412\ : InMux
    port map (
            O => \N__42496\,
            I => \N__42489\
        );

    \I__9411\ : InMux
    port map (
            O => \N__42493\,
            I => \N__42484\
        );

    \I__9410\ : InMux
    port map (
            O => \N__42492\,
            I => \N__42484\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__42489\,
            I => \N__42481\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__42484\,
            I => \N__42478\
        );

    \I__9407\ : Span4Mux_h
    port map (
            O => \N__42481\,
            I => \N__42474\
        );

    \I__9406\ : Span12Mux_v
    port map (
            O => \N__42478\,
            I => \N__42471\
        );

    \I__9405\ : InMux
    port map (
            O => \N__42477\,
            I => \N__42468\
        );

    \I__9404\ : Odrv4
    port map (
            O => \N__42474\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9403\ : Odrv12
    port map (
            O => \N__42471\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__42468\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9401\ : InMux
    port map (
            O => \N__42461\,
            I => \N__42458\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__42458\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__9399\ : CascadeMux
    port map (
            O => \N__42455\,
            I => \N__42452\
        );

    \I__9398\ : InMux
    port map (
            O => \N__42452\,
            I => \N__42449\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__42449\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__9396\ : InMux
    port map (
            O => \N__42446\,
            I => \N__42443\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__42443\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__9394\ : InMux
    port map (
            O => \N__42440\,
            I => \N__42436\
        );

    \I__9393\ : InMux
    port map (
            O => \N__42439\,
            I => \N__42433\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__42436\,
            I => \N__42430\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__42433\,
            I => \current_shift_inst.un4_control_input_0_31\
        );

    \I__9390\ : Odrv12
    port map (
            O => \N__42430\,
            I => \current_shift_inst.un4_control_input_0_31\
        );

    \I__9389\ : CascadeMux
    port map (
            O => \N__42425\,
            I => \N__42422\
        );

    \I__9388\ : InMux
    port map (
            O => \N__42422\,
            I => \N__42419\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__42419\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__9386\ : InMux
    port map (
            O => \N__42416\,
            I => \N__42413\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__42413\,
            I => \N__42410\
        );

    \I__9384\ : Odrv4
    port map (
            O => \N__42410\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__9383\ : CascadeMux
    port map (
            O => \N__42407\,
            I => \N__42404\
        );

    \I__9382\ : InMux
    port map (
            O => \N__42404\,
            I => \N__42401\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__42401\,
            I => \N__42398\
        );

    \I__9380\ : Odrv12
    port map (
            O => \N__42398\,
            I => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\
        );

    \I__9379\ : InMux
    port map (
            O => \N__42395\,
            I => \N__42392\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__42392\,
            I => \N__42389\
        );

    \I__9377\ : Odrv4
    port map (
            O => \N__42389\,
            I => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\
        );

    \I__9376\ : InMux
    port map (
            O => \N__42386\,
            I => \N__42383\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__42383\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__9374\ : InMux
    port map (
            O => \N__42380\,
            I => \N__42377\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__42377\,
            I => \N__42374\
        );

    \I__9372\ : Odrv12
    port map (
            O => \N__42374\,
            I => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\
        );

    \I__9371\ : InMux
    port map (
            O => \N__42371\,
            I => \N__42368\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__42368\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__9369\ : InMux
    port map (
            O => \N__42365\,
            I => \N__42362\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__42362\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__9367\ : CascadeMux
    port map (
            O => \N__42359\,
            I => \N__42356\
        );

    \I__9366\ : InMux
    port map (
            O => \N__42356\,
            I => \N__42353\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__42353\,
            I => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\
        );

    \I__9364\ : CascadeMux
    port map (
            O => \N__42350\,
            I => \N__42347\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42347\,
            I => \N__42344\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__42344\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__9361\ : CascadeMux
    port map (
            O => \N__42341\,
            I => \N__42338\
        );

    \I__9360\ : InMux
    port map (
            O => \N__42338\,
            I => \N__42335\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__42335\,
            I => \N__42332\
        );

    \I__9358\ : Odrv4
    port map (
            O => \N__42332\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__9357\ : InMux
    port map (
            O => \N__42329\,
            I => \N__42326\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__42326\,
            I => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\
        );

    \I__9355\ : InMux
    port map (
            O => \N__42323\,
            I => \N__42320\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__42320\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__9353\ : CascadeMux
    port map (
            O => \N__42317\,
            I => \N__42314\
        );

    \I__9352\ : InMux
    port map (
            O => \N__42314\,
            I => \N__42311\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__42311\,
            I => \N__42308\
        );

    \I__9350\ : Odrv12
    port map (
            O => \N__42308\,
            I => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\
        );

    \I__9349\ : CascadeMux
    port map (
            O => \N__42305\,
            I => \N__42302\
        );

    \I__9348\ : InMux
    port map (
            O => \N__42302\,
            I => \N__42299\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__42299\,
            I => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\
        );

    \I__9346\ : CascadeMux
    port map (
            O => \N__42296\,
            I => \N__42293\
        );

    \I__9345\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42290\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__42290\,
            I => \N__42287\
        );

    \I__9343\ : Odrv4
    port map (
            O => \N__42287\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__9342\ : InMux
    port map (
            O => \N__42284\,
            I => \N__42281\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__42281\,
            I => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\
        );

    \I__9340\ : InMux
    port map (
            O => \N__42278\,
            I => \N__42275\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__42275\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__9338\ : InMux
    port map (
            O => \N__42272\,
            I => \bfn_16_17_0_\
        );

    \I__9337\ : InMux
    port map (
            O => \N__42269\,
            I => \N__42266\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__42266\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__9335\ : InMux
    port map (
            O => \N__42263\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__9334\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42257\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__42257\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__9332\ : InMux
    port map (
            O => \N__42254\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__9331\ : CascadeMux
    port map (
            O => \N__42251\,
            I => \N__42248\
        );

    \I__9330\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42245\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__42245\,
            I => \N__42242\
        );

    \I__9328\ : Span4Mux_v
    port map (
            O => \N__42242\,
            I => \N__42239\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__42239\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__9326\ : InMux
    port map (
            O => \N__42236\,
            I => \N__42233\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__42233\,
            I => \N__42230\
        );

    \I__9324\ : Odrv4
    port map (
            O => \N__42230\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__9323\ : InMux
    port map (
            O => \N__42227\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__9322\ : InMux
    port map (
            O => \N__42224\,
            I => \N__42221\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__42221\,
            I => \N__42218\
        );

    \I__9320\ : Odrv4
    port map (
            O => \N__42218\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42215\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__9318\ : InMux
    port map (
            O => \N__42212\,
            I => \N__42209\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__42209\,
            I => \N__42206\
        );

    \I__9316\ : Odrv4
    port map (
            O => \N__42206\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__9315\ : InMux
    port map (
            O => \N__42203\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__9314\ : InMux
    port map (
            O => \N__42200\,
            I => \N__42197\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__42197\,
            I => \N__42194\
        );

    \I__9312\ : Odrv4
    port map (
            O => \N__42194\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__9311\ : InMux
    port map (
            O => \N__42191\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__9310\ : InMux
    port map (
            O => \N__42188\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__9309\ : InMux
    port map (
            O => \N__42185\,
            I => \N__42182\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__42182\,
            I => \N__42179\
        );

    \I__9307\ : Odrv4
    port map (
            O => \N__42179\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__9306\ : CascadeMux
    port map (
            O => \N__42176\,
            I => \N__42173\
        );

    \I__9305\ : InMux
    port map (
            O => \N__42173\,
            I => \N__42170\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__42170\,
            I => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\
        );

    \I__9303\ : InMux
    port map (
            O => \N__42167\,
            I => \N__42164\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__42164\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__9301\ : InMux
    port map (
            O => \N__42161\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__9300\ : InMux
    port map (
            O => \N__42158\,
            I => \N__42155\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__42155\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__9298\ : InMux
    port map (
            O => \N__42152\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__9297\ : InMux
    port map (
            O => \N__42149\,
            I => \N__42146\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__42146\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__9295\ : InMux
    port map (
            O => \N__42143\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__9294\ : InMux
    port map (
            O => \N__42140\,
            I => \N__42137\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__42137\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__9292\ : InMux
    port map (
            O => \N__42134\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__9291\ : CascadeMux
    port map (
            O => \N__42131\,
            I => \N__42128\
        );

    \I__9290\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42125\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__42125\,
            I => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\
        );

    \I__9288\ : InMux
    port map (
            O => \N__42122\,
            I => \N__42119\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__42119\,
            I => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\
        );

    \I__9286\ : InMux
    port map (
            O => \N__42116\,
            I => \N__42113\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__42113\,
            I => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\
        );

    \I__9284\ : InMux
    port map (
            O => \N__42110\,
            I => \N__42106\
        );

    \I__9283\ : InMux
    port map (
            O => \N__42109\,
            I => \N__42103\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__42106\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__42103\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9280\ : InMux
    port map (
            O => \N__42098\,
            I => \N__42095\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__42095\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__9278\ : InMux
    port map (
            O => \N__42092\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__9277\ : InMux
    port map (
            O => \N__42089\,
            I => \N__42085\
        );

    \I__9276\ : InMux
    port map (
            O => \N__42088\,
            I => \N__42082\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__42085\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__42082\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9273\ : InMux
    port map (
            O => \N__42077\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__9272\ : InMux
    port map (
            O => \N__42074\,
            I => \N__42071\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__42071\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__9270\ : InMux
    port map (
            O => \N__42068\,
            I => \N__42065\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__42065\,
            I => \N__42061\
        );

    \I__9268\ : InMux
    port map (
            O => \N__42064\,
            I => \N__42058\
        );

    \I__9267\ : Span4Mux_h
    port map (
            O => \N__42061\,
            I => \N__42055\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__42058\,
            I => \N__42052\
        );

    \I__9265\ : Span4Mux_v
    port map (
            O => \N__42055\,
            I => \N__42049\
        );

    \I__9264\ : Odrv12
    port map (
            O => \N__42052\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__9263\ : Odrv4
    port map (
            O => \N__42049\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__9262\ : CascadeMux
    port map (
            O => \N__42044\,
            I => \N__42040\
        );

    \I__9261\ : CascadeMux
    port map (
            O => \N__42043\,
            I => \N__42037\
        );

    \I__9260\ : InMux
    port map (
            O => \N__42040\,
            I => \N__42034\
        );

    \I__9259\ : InMux
    port map (
            O => \N__42037\,
            I => \N__42031\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__42034\,
            I => \N__42028\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__42031\,
            I => \N__42025\
        );

    \I__9256\ : Span12Mux_s11_h
    port map (
            O => \N__42028\,
            I => \N__42022\
        );

    \I__9255\ : Span4Mux_v
    port map (
            O => \N__42025\,
            I => \N__42019\
        );

    \I__9254\ : Odrv12
    port map (
            O => \N__42022\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__9253\ : Odrv4
    port map (
            O => \N__42019\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__9252\ : InMux
    port map (
            O => \N__42014\,
            I => \N__42011\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__42011\,
            I => \N__42008\
        );

    \I__9250\ : Span4Mux_h
    port map (
            O => \N__42008\,
            I => \N__42005\
        );

    \I__9249\ : Span4Mux_h
    port map (
            O => \N__42005\,
            I => \N__42002\
        );

    \I__9248\ : Odrv4
    port map (
            O => \N__42002\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__9247\ : InMux
    port map (
            O => \N__41999\,
            I => \N__41996\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__41996\,
            I => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\
        );

    \I__9245\ : InMux
    port map (
            O => \N__41993\,
            I => \N__41990\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__41990\,
            I => \N__41987\
        );

    \I__9243\ : Span4Mux_h
    port map (
            O => \N__41987\,
            I => \N__41983\
        );

    \I__9242\ : InMux
    port map (
            O => \N__41986\,
            I => \N__41980\
        );

    \I__9241\ : Odrv4
    port map (
            O => \N__41983\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__41980\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__9239\ : InMux
    port map (
            O => \N__41975\,
            I => \N__41972\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__41972\,
            I => \N__41969\
        );

    \I__9237\ : Span4Mux_v
    port map (
            O => \N__41969\,
            I => \N__41966\
        );

    \I__9236\ : Odrv4
    port map (
            O => \N__41966\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__9235\ : InMux
    port map (
            O => \N__41963\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__9234\ : InMux
    port map (
            O => \N__41960\,
            I => \N__41957\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__41957\,
            I => \N__41954\
        );

    \I__9232\ : Span4Mux_h
    port map (
            O => \N__41954\,
            I => \N__41950\
        );

    \I__9231\ : InMux
    port map (
            O => \N__41953\,
            I => \N__41947\
        );

    \I__9230\ : Odrv4
    port map (
            O => \N__41950\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__41947\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__9228\ : InMux
    port map (
            O => \N__41942\,
            I => \N__41939\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__41939\,
            I => \N__41936\
        );

    \I__9226\ : Span4Mux_h
    port map (
            O => \N__41936\,
            I => \N__41933\
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__41933\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__9224\ : InMux
    port map (
            O => \N__41930\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__9223\ : InMux
    port map (
            O => \N__41927\,
            I => \N__41924\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__41924\,
            I => \N__41921\
        );

    \I__9221\ : Span4Mux_v
    port map (
            O => \N__41921\,
            I => \N__41917\
        );

    \I__9220\ : InMux
    port map (
            O => \N__41920\,
            I => \N__41914\
        );

    \I__9219\ : Odrv4
    port map (
            O => \N__41917\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__41914\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__9217\ : InMux
    port map (
            O => \N__41909\,
            I => \N__41906\
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__41906\,
            I => \N__41903\
        );

    \I__9215\ : Span4Mux_h
    port map (
            O => \N__41903\,
            I => \N__41900\
        );

    \I__9214\ : Odrv4
    port map (
            O => \N__41900\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__9213\ : InMux
    port map (
            O => \N__41897\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__9212\ : InMux
    port map (
            O => \N__41894\,
            I => \N__41891\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__41891\,
            I => \N__41888\
        );

    \I__9210\ : Span4Mux_v
    port map (
            O => \N__41888\,
            I => \N__41884\
        );

    \I__9209\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41881\
        );

    \I__9208\ : Odrv4
    port map (
            O => \N__41884\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__41881\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__9206\ : InMux
    port map (
            O => \N__41876\,
            I => \N__41873\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41873\,
            I => \N__41870\
        );

    \I__9204\ : Span4Mux_h
    port map (
            O => \N__41870\,
            I => \N__41867\
        );

    \I__9203\ : Odrv4
    port map (
            O => \N__41867\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__9202\ : InMux
    port map (
            O => \N__41864\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__9201\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41858\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__41858\,
            I => \N__41855\
        );

    \I__9199\ : Span4Mux_h
    port map (
            O => \N__41855\,
            I => \N__41851\
        );

    \I__9198\ : InMux
    port map (
            O => \N__41854\,
            I => \N__41848\
        );

    \I__9197\ : Odrv4
    port map (
            O => \N__41851\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__41848\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41843\,
            I => \N__41840\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__41840\,
            I => \N__41837\
        );

    \I__9193\ : Span4Mux_h
    port map (
            O => \N__41837\,
            I => \N__41834\
        );

    \I__9192\ : Odrv4
    port map (
            O => \N__41834\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__9191\ : InMux
    port map (
            O => \N__41831\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__9190\ : InMux
    port map (
            O => \N__41828\,
            I => \N__41825\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__41825\,
            I => \N__41822\
        );

    \I__9188\ : Span4Mux_h
    port map (
            O => \N__41822\,
            I => \N__41818\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41821\,
            I => \N__41815\
        );

    \I__9186\ : Odrv4
    port map (
            O => \N__41818\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__41815\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9184\ : InMux
    port map (
            O => \N__41810\,
            I => \N__41807\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__41807\,
            I => \N__41804\
        );

    \I__9182\ : Span4Mux_h
    port map (
            O => \N__41804\,
            I => \N__41801\
        );

    \I__9181\ : Odrv4
    port map (
            O => \N__41801\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__9180\ : InMux
    port map (
            O => \N__41798\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__9179\ : InMux
    port map (
            O => \N__41795\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__9178\ : InMux
    port map (
            O => \N__41792\,
            I => \N__41788\
        );

    \I__9177\ : InMux
    port map (
            O => \N__41791\,
            I => \N__41785\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__41788\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__41785\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9174\ : InMux
    port map (
            O => \N__41780\,
            I => \N__41777\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__41777\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__9172\ : InMux
    port map (
            O => \N__41774\,
            I => \bfn_16_13_0_\
        );

    \I__9171\ : InMux
    port map (
            O => \N__41771\,
            I => \N__41768\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__41768\,
            I => \N__41765\
        );

    \I__9169\ : Odrv4
    port map (
            O => \N__41765\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__9168\ : InMux
    port map (
            O => \N__41762\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__9167\ : InMux
    port map (
            O => \N__41759\,
            I => \N__41756\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__41756\,
            I => \N__41753\
        );

    \I__9165\ : Span4Mux_h
    port map (
            O => \N__41753\,
            I => \N__41750\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__41750\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\
        );

    \I__9163\ : CascadeMux
    port map (
            O => \N__41747\,
            I => \N__41744\
        );

    \I__9162\ : InMux
    port map (
            O => \N__41744\,
            I => \N__41740\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41743\,
            I => \N__41737\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__41740\,
            I => \N__41734\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__41737\,
            I => \N__41731\
        );

    \I__9158\ : Odrv4
    port map (
            O => \N__41734\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__9157\ : Odrv4
    port map (
            O => \N__41731\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__9156\ : InMux
    port map (
            O => \N__41726\,
            I => \N__41723\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__41723\,
            I => \N__41720\
        );

    \I__9154\ : Odrv4
    port map (
            O => \N__41720\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__9153\ : InMux
    port map (
            O => \N__41717\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__9152\ : InMux
    port map (
            O => \N__41714\,
            I => \N__41710\
        );

    \I__9151\ : InMux
    port map (
            O => \N__41713\,
            I => \N__41707\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__41710\,
            I => \N__41704\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__41707\,
            I => \N__41701\
        );

    \I__9148\ : Odrv4
    port map (
            O => \N__41704\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__9147\ : Odrv4
    port map (
            O => \N__41701\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__9146\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41693\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__41693\,
            I => \N__41690\
        );

    \I__9144\ : Odrv4
    port map (
            O => \N__41690\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__9143\ : InMux
    port map (
            O => \N__41687\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__9142\ : InMux
    port map (
            O => \N__41684\,
            I => \N__41680\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41683\,
            I => \N__41677\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__41680\,
            I => \N__41674\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__41677\,
            I => \N__41671\
        );

    \I__9138\ : Odrv4
    port map (
            O => \N__41674\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__9137\ : Odrv12
    port map (
            O => \N__41671\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__9136\ : InMux
    port map (
            O => \N__41666\,
            I => \N__41663\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__41663\,
            I => \N__41660\
        );

    \I__9134\ : Odrv4
    port map (
            O => \N__41660\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__9133\ : InMux
    port map (
            O => \N__41657\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41654\,
            I => \N__41651\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__41651\,
            I => \N__41647\
        );

    \I__9130\ : InMux
    port map (
            O => \N__41650\,
            I => \N__41644\
        );

    \I__9129\ : Span4Mux_v
    port map (
            O => \N__41647\,
            I => \N__41639\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41644\,
            I => \N__41639\
        );

    \I__9127\ : Span4Mux_h
    port map (
            O => \N__41639\,
            I => \N__41636\
        );

    \I__9126\ : Odrv4
    port map (
            O => \N__41636\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41633\,
            I => \N__41630\
        );

    \I__9124\ : LocalMux
    port map (
            O => \N__41630\,
            I => \N__41627\
        );

    \I__9123\ : Odrv4
    port map (
            O => \N__41627\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__9122\ : InMux
    port map (
            O => \N__41624\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__9121\ : InMux
    port map (
            O => \N__41621\,
            I => \N__41618\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__41618\,
            I => \N__41614\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41617\,
            I => \N__41611\
        );

    \I__9118\ : Span4Mux_v
    port map (
            O => \N__41614\,
            I => \N__41608\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41611\,
            I => \N__41605\
        );

    \I__9116\ : Odrv4
    port map (
            O => \N__41608\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9115\ : Odrv4
    port map (
            O => \N__41605\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41597\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__41597\,
            I => \N__41594\
        );

    \I__9112\ : Span4Mux_h
    port map (
            O => \N__41594\,
            I => \N__41591\
        );

    \I__9111\ : Odrv4
    port map (
            O => \N__41591\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__9110\ : InMux
    port map (
            O => \N__41588\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41585\,
            I => \N__41581\
        );

    \I__9108\ : InMux
    port map (
            O => \N__41584\,
            I => \N__41578\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__41581\,
            I => \N__41575\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__41578\,
            I => \N__41572\
        );

    \I__9105\ : Span4Mux_v
    port map (
            O => \N__41575\,
            I => \N__41569\
        );

    \I__9104\ : Span4Mux_h
    port map (
            O => \N__41572\,
            I => \N__41566\
        );

    \I__9103\ : Odrv4
    port map (
            O => \N__41569\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9102\ : Odrv4
    port map (
            O => \N__41566\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9101\ : InMux
    port map (
            O => \N__41561\,
            I => \N__41558\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__41558\,
            I => \N__41555\
        );

    \I__9099\ : Span4Mux_h
    port map (
            O => \N__41555\,
            I => \N__41552\
        );

    \I__9098\ : Odrv4
    port map (
            O => \N__41552\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41549\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41546\,
            I => \N__41543\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__41543\,
            I => \N__41539\
        );

    \I__9094\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41536\
        );

    \I__9093\ : Odrv4
    port map (
            O => \N__41539\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__41536\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41531\,
            I => \N__41528\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__41528\,
            I => \N__41525\
        );

    \I__9089\ : Odrv4
    port map (
            O => \N__41525\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__9088\ : InMux
    port map (
            O => \N__41522\,
            I => \bfn_16_12_0_\
        );

    \I__9087\ : InMux
    port map (
            O => \N__41519\,
            I => \N__41516\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__41516\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__9085\ : InMux
    port map (
            O => \N__41513\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41510\,
            I => \N__41507\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__41507\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9082\ : InMux
    port map (
            O => \N__41504\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__9081\ : CascadeMux
    port map (
            O => \N__41501\,
            I => \N__41498\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41498\,
            I => \N__41495\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__41495\,
            I => \N__41492\
        );

    \I__9078\ : Odrv4
    port map (
            O => \N__41492\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41489\,
            I => \bfn_16_10_0_\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41486\,
            I => \N__41483\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__41483\,
            I => \N__41480\
        );

    \I__9074\ : Span4Mux_h
    port map (
            O => \N__41480\,
            I => \N__41477\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__41477\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__9072\ : InMux
    port map (
            O => \N__41474\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__9071\ : InMux
    port map (
            O => \N__41471\,
            I => \N__41468\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__41468\,
            I => \N__41465\
        );

    \I__9069\ : Span4Mux_h
    port map (
            O => \N__41465\,
            I => \N__41462\
        );

    \I__9068\ : Odrv4
    port map (
            O => \N__41462\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9067\ : InMux
    port map (
            O => \N__41459\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__9066\ : CascadeMux
    port map (
            O => \N__41456\,
            I => \N__41453\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41453\,
            I => \N__41450\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__41450\,
            I => \N__41447\
        );

    \I__9063\ : Span4Mux_h
    port map (
            O => \N__41447\,
            I => \N__41444\
        );

    \I__9062\ : Odrv4
    port map (
            O => \N__41444\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__9061\ : InMux
    port map (
            O => \N__41441\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41438\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__9059\ : CascadeMux
    port map (
            O => \N__41435\,
            I => \N__41430\
        );

    \I__9058\ : InMux
    port map (
            O => \N__41434\,
            I => \N__41418\
        );

    \I__9057\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41418\
        );

    \I__9056\ : InMux
    port map (
            O => \N__41430\,
            I => \N__41418\
        );

    \I__9055\ : InMux
    port map (
            O => \N__41429\,
            I => \N__41418\
        );

    \I__9054\ : CascadeMux
    port map (
            O => \N__41428\,
            I => \N__41414\
        );

    \I__9053\ : CascadeMux
    port map (
            O => \N__41427\,
            I => \N__41411\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__41418\,
            I => \N__41402\
        );

    \I__9051\ : CascadeMux
    port map (
            O => \N__41417\,
            I => \N__41399\
        );

    \I__9050\ : InMux
    port map (
            O => \N__41414\,
            I => \N__41396\
        );

    \I__9049\ : InMux
    port map (
            O => \N__41411\,
            I => \N__41383\
        );

    \I__9048\ : InMux
    port map (
            O => \N__41410\,
            I => \N__41383\
        );

    \I__9047\ : InMux
    port map (
            O => \N__41409\,
            I => \N__41383\
        );

    \I__9046\ : InMux
    port map (
            O => \N__41408\,
            I => \N__41383\
        );

    \I__9045\ : InMux
    port map (
            O => \N__41407\,
            I => \N__41383\
        );

    \I__9044\ : InMux
    port map (
            O => \N__41406\,
            I => \N__41383\
        );

    \I__9043\ : CascadeMux
    port map (
            O => \N__41405\,
            I => \N__41380\
        );

    \I__9042\ : Span4Mux_v
    port map (
            O => \N__41402\,
            I => \N__41377\
        );

    \I__9041\ : InMux
    port map (
            O => \N__41399\,
            I => \N__41374\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__41396\,
            I => \N__41371\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__41383\,
            I => \N__41368\
        );

    \I__9038\ : InMux
    port map (
            O => \N__41380\,
            I => \N__41365\
        );

    \I__9037\ : Span4Mux_h
    port map (
            O => \N__41377\,
            I => \N__41360\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__41374\,
            I => \N__41360\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__41371\,
            I => \N__41353\
        );

    \I__9034\ : Span4Mux_h
    port map (
            O => \N__41368\,
            I => \N__41353\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__41365\,
            I => \N__41353\
        );

    \I__9032\ : Sp12to4
    port map (
            O => \N__41360\,
            I => \N__41350\
        );

    \I__9031\ : Span4Mux_v
    port map (
            O => \N__41353\,
            I => \N__41347\
        );

    \I__9030\ : Odrv12
    port map (
            O => \N__41350\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__41347\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__9028\ : InMux
    port map (
            O => \N__41342\,
            I => \N__41339\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__41339\,
            I => \N__41336\
        );

    \I__9026\ : Span4Mux_h
    port map (
            O => \N__41336\,
            I => \N__41333\
        );

    \I__9025\ : Odrv4
    port map (
            O => \N__41333\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__9024\ : CascadeMux
    port map (
            O => \N__41330\,
            I => \N__41326\
        );

    \I__9023\ : InMux
    port map (
            O => \N__41329\,
            I => \N__41323\
        );

    \I__9022\ : InMux
    port map (
            O => \N__41326\,
            I => \N__41320\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__41323\,
            I => \N__41314\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__41320\,
            I => \N__41314\
        );

    \I__9019\ : InMux
    port map (
            O => \N__41319\,
            I => \N__41311\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__41314\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__41311\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__9016\ : InMux
    port map (
            O => \N__41306\,
            I => \N__41302\
        );

    \I__9015\ : InMux
    port map (
            O => \N__41305\,
            I => \N__41299\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__41302\,
            I => \N__41296\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41299\,
            I => \N__41293\
        );

    \I__9012\ : Odrv4
    port map (
            O => \N__41296\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__9011\ : Odrv4
    port map (
            O => \N__41293\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__9010\ : InMux
    port map (
            O => \N__41288\,
            I => \N__41285\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__41285\,
            I => \N__41282\
        );

    \I__9008\ : Span4Mux_h
    port map (
            O => \N__41282\,
            I => \N__41277\
        );

    \I__9007\ : InMux
    port map (
            O => \N__41281\,
            I => \N__41272\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41280\,
            I => \N__41272\
        );

    \I__9005\ : Span4Mux_h
    port map (
            O => \N__41277\,
            I => \N__41267\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__41272\,
            I => \N__41267\
        );

    \I__9003\ : Odrv4
    port map (
            O => \N__41267\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__9002\ : InMux
    port map (
            O => \N__41264\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__9001\ : InMux
    port map (
            O => \N__41261\,
            I => \N__41258\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41258\,
            I => \N__41253\
        );

    \I__8999\ : InMux
    port map (
            O => \N__41257\,
            I => \N__41248\
        );

    \I__8998\ : InMux
    port map (
            O => \N__41256\,
            I => \N__41248\
        );

    \I__8997\ : Span4Mux_v
    port map (
            O => \N__41253\,
            I => \N__41245\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__41248\,
            I => \N__41242\
        );

    \I__8995\ : Odrv4
    port map (
            O => \N__41245\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__8994\ : Odrv4
    port map (
            O => \N__41242\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__8993\ : InMux
    port map (
            O => \N__41237\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__8992\ : InMux
    port map (
            O => \N__41234\,
            I => \N__41229\
        );

    \I__8991\ : CascadeMux
    port map (
            O => \N__41233\,
            I => \N__41226\
        );

    \I__8990\ : CascadeMux
    port map (
            O => \N__41232\,
            I => \N__41223\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__41229\,
            I => \N__41220\
        );

    \I__8988\ : InMux
    port map (
            O => \N__41226\,
            I => \N__41215\
        );

    \I__8987\ : InMux
    port map (
            O => \N__41223\,
            I => \N__41215\
        );

    \I__8986\ : Span12Mux_h
    port map (
            O => \N__41220\,
            I => \N__41212\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__41215\,
            I => \N__41209\
        );

    \I__8984\ : Odrv12
    port map (
            O => \N__41212\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__8983\ : Odrv4
    port map (
            O => \N__41209\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__8982\ : InMux
    port map (
            O => \N__41204\,
            I => \bfn_16_9_0_\
        );

    \I__8981\ : InMux
    port map (
            O => \N__41201\,
            I => \N__41198\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__41198\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__8979\ : InMux
    port map (
            O => \N__41195\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__8978\ : InMux
    port map (
            O => \N__41192\,
            I => \N__41189\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__41189\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__8976\ : InMux
    port map (
            O => \N__41186\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8975\ : InMux
    port map (
            O => \N__41183\,
            I => \N__41180\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__41180\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__8973\ : InMux
    port map (
            O => \N__41177\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8972\ : CascadeMux
    port map (
            O => \N__41174\,
            I => \N__41171\
        );

    \I__8971\ : InMux
    port map (
            O => \N__41171\,
            I => \N__41168\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__41168\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__8969\ : InMux
    port map (
            O => \N__41165\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8968\ : InMux
    port map (
            O => \N__41162\,
            I => \N__41159\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__41159\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__8966\ : InMux
    port map (
            O => \N__41156\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8965\ : InMux
    port map (
            O => \N__41153\,
            I => \N__41150\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__41150\,
            I => \N__41146\
        );

    \I__8963\ : InMux
    port map (
            O => \N__41149\,
            I => \N__41143\
        );

    \I__8962\ : Span12Mux_v
    port map (
            O => \N__41146\,
            I => \N__41140\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__41143\,
            I => \N__41137\
        );

    \I__8960\ : Odrv12
    port map (
            O => \N__41140\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__8959\ : Odrv12
    port map (
            O => \N__41137\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__8958\ : InMux
    port map (
            O => \N__41132\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__8957\ : InMux
    port map (
            O => \N__41129\,
            I => \N__41125\
        );

    \I__8956\ : InMux
    port map (
            O => \N__41128\,
            I => \N__41122\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__41125\,
            I => \N__41116\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__41122\,
            I => \N__41116\
        );

    \I__8953\ : InMux
    port map (
            O => \N__41121\,
            I => \N__41113\
        );

    \I__8952\ : Span4Mux_h
    port map (
            O => \N__41116\,
            I => \N__41108\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__41113\,
            I => \N__41105\
        );

    \I__8950\ : InMux
    port map (
            O => \N__41112\,
            I => \N__41102\
        );

    \I__8949\ : InMux
    port map (
            O => \N__41111\,
            I => \N__41099\
        );

    \I__8948\ : Span4Mux_h
    port map (
            O => \N__41108\,
            I => \N__41096\
        );

    \I__8947\ : Span4Mux_v
    port map (
            O => \N__41105\,
            I => \N__41093\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__41102\,
            I => \N__41088\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__41099\,
            I => \N__41088\
        );

    \I__8944\ : Odrv4
    port map (
            O => \N__41096\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__8943\ : Odrv4
    port map (
            O => \N__41093\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__8942\ : Odrv12
    port map (
            O => \N__41088\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__8941\ : InMux
    port map (
            O => \N__41081\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__8940\ : InMux
    port map (
            O => \N__41078\,
            I => \N__41075\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__41075\,
            I => \N__41071\
        );

    \I__8938\ : InMux
    port map (
            O => \N__41074\,
            I => \N__41068\
        );

    \I__8937\ : Span4Mux_v
    port map (
            O => \N__41071\,
            I => \N__41065\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__41068\,
            I => \N__41062\
        );

    \I__8935\ : Odrv4
    port map (
            O => \N__41065\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__8934\ : Odrv12
    port map (
            O => \N__41062\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__8933\ : InMux
    port map (
            O => \N__41057\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__8932\ : InMux
    port map (
            O => \N__41054\,
            I => \N__41050\
        );

    \I__8931\ : InMux
    port map (
            O => \N__41053\,
            I => \N__41047\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__41050\,
            I => \N__41042\
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__41047\,
            I => \N__41042\
        );

    \I__8928\ : Span12Mux_s7_v
    port map (
            O => \N__41042\,
            I => \N__41039\
        );

    \I__8927\ : Odrv12
    port map (
            O => \N__41039\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__8926\ : InMux
    port map (
            O => \N__41036\,
            I => \bfn_16_8_0_\
        );

    \I__8925\ : InMux
    port map (
            O => \N__41033\,
            I => \N__41029\
        );

    \I__8924\ : InMux
    port map (
            O => \N__41032\,
            I => \N__41026\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__41029\,
            I => \N__41021\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__41026\,
            I => \N__41021\
        );

    \I__8921\ : Span4Mux_v
    port map (
            O => \N__41021\,
            I => \N__41018\
        );

    \I__8920\ : Span4Mux_h
    port map (
            O => \N__41018\,
            I => \N__41015\
        );

    \I__8919\ : Odrv4
    port map (
            O => \N__41015\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__8918\ : InMux
    port map (
            O => \N__41012\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__8917\ : CascadeMux
    port map (
            O => \N__41009\,
            I => \N__41005\
        );

    \I__8916\ : InMux
    port map (
            O => \N__41008\,
            I => \N__41002\
        );

    \I__8915\ : InMux
    port map (
            O => \N__41005\,
            I => \N__40999\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__41002\,
            I => \N__40994\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__40999\,
            I => \N__40994\
        );

    \I__8912\ : Span4Mux_v
    port map (
            O => \N__40994\,
            I => \N__40991\
        );

    \I__8911\ : Odrv4
    port map (
            O => \N__40991\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__8910\ : InMux
    port map (
            O => \N__40988\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8909\ : InMux
    port map (
            O => \N__40985\,
            I => \N__40980\
        );

    \I__8908\ : InMux
    port map (
            O => \N__40984\,
            I => \N__40977\
        );

    \I__8907\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40972\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__40980\,
            I => \N__40967\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__40977\,
            I => \N__40967\
        );

    \I__8904\ : InMux
    port map (
            O => \N__40976\,
            I => \N__40964\
        );

    \I__8903\ : InMux
    port map (
            O => \N__40975\,
            I => \N__40961\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__40972\,
            I => \N__40958\
        );

    \I__8901\ : Span4Mux_v
    port map (
            O => \N__40967\,
            I => \N__40951\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__40964\,
            I => \N__40951\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__40961\,
            I => \N__40951\
        );

    \I__8898\ : Span4Mux_v
    port map (
            O => \N__40958\,
            I => \N__40948\
        );

    \I__8897\ : Span4Mux_h
    port map (
            O => \N__40951\,
            I => \N__40945\
        );

    \I__8896\ : Odrv4
    port map (
            O => \N__40948\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__8895\ : Odrv4
    port map (
            O => \N__40945\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__8894\ : InMux
    port map (
            O => \N__40940\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__8893\ : InMux
    port map (
            O => \N__40937\,
            I => \N__40929\
        );

    \I__8892\ : InMux
    port map (
            O => \N__40936\,
            I => \N__40929\
        );

    \I__8891\ : InMux
    port map (
            O => \N__40935\,
            I => \N__40925\
        );

    \I__8890\ : CascadeMux
    port map (
            O => \N__40934\,
            I => \N__40921\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__40929\,
            I => \N__40918\
        );

    \I__8888\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40915\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__40925\,
            I => \N__40912\
        );

    \I__8886\ : InMux
    port map (
            O => \N__40924\,
            I => \N__40907\
        );

    \I__8885\ : InMux
    port map (
            O => \N__40921\,
            I => \N__40907\
        );

    \I__8884\ : Span4Mux_h
    port map (
            O => \N__40918\,
            I => \N__40904\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__40915\,
            I => \N__40901\
        );

    \I__8882\ : Span4Mux_h
    port map (
            O => \N__40912\,
            I => \N__40896\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__40907\,
            I => \N__40896\
        );

    \I__8880\ : Span4Mux_h
    port map (
            O => \N__40904\,
            I => \N__40893\
        );

    \I__8879\ : Span4Mux_v
    port map (
            O => \N__40901\,
            I => \N__40888\
        );

    \I__8878\ : Span4Mux_v
    port map (
            O => \N__40896\,
            I => \N__40888\
        );

    \I__8877\ : Odrv4
    port map (
            O => \N__40893\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8876\ : Odrv4
    port map (
            O => \N__40888\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8875\ : InMux
    port map (
            O => \N__40883\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__8874\ : InMux
    port map (
            O => \N__40880\,
            I => \N__40877\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__40877\,
            I => \N__40874\
        );

    \I__8872\ : Span4Mux_v
    port map (
            O => \N__40874\,
            I => \N__40869\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40873\,
            I => \N__40866\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40872\,
            I => \N__40863\
        );

    \I__8869\ : Span4Mux_h
    port map (
            O => \N__40869\,
            I => \N__40856\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__40866\,
            I => \N__40856\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__40863\,
            I => \N__40856\
        );

    \I__8866\ : Odrv4
    port map (
            O => \N__40856\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__8865\ : InMux
    port map (
            O => \N__40853\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__8864\ : CascadeMux
    port map (
            O => \N__40850\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\
        );

    \I__8863\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40844\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__40844\,
            I => \N__40841\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__40841\,
            I => \N__40838\
        );

    \I__8860\ : Odrv4
    port map (
            O => \N__40838\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\
        );

    \I__8859\ : CascadeMux
    port map (
            O => \N__40835\,
            I => \N__40830\
        );

    \I__8858\ : InMux
    port map (
            O => \N__40834\,
            I => \N__40826\
        );

    \I__8857\ : InMux
    port map (
            O => \N__40833\,
            I => \N__40823\
        );

    \I__8856\ : InMux
    port map (
            O => \N__40830\,
            I => \N__40820\
        );

    \I__8855\ : InMux
    port map (
            O => \N__40829\,
            I => \N__40817\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__40826\,
            I => \N__40814\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__40823\,
            I => \N__40811\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__40820\,
            I => \N__40808\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__40817\,
            I => \N__40805\
        );

    \I__8850\ : Span4Mux_v
    port map (
            O => \N__40814\,
            I => \N__40800\
        );

    \I__8849\ : Span4Mux_v
    port map (
            O => \N__40811\,
            I => \N__40800\
        );

    \I__8848\ : Odrv12
    port map (
            O => \N__40808\,
            I => \delay_measurement_inst.N_265\
        );

    \I__8847\ : Odrv4
    port map (
            O => \N__40805\,
            I => \delay_measurement_inst.N_265\
        );

    \I__8846\ : Odrv4
    port map (
            O => \N__40800\,
            I => \delay_measurement_inst.N_265\
        );

    \I__8845\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40790\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__40790\,
            I => \N__40787\
        );

    \I__8843\ : Span4Mux_h
    port map (
            O => \N__40787\,
            I => \N__40783\
        );

    \I__8842\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40780\
        );

    \I__8841\ : Odrv4
    port map (
            O => \N__40783\,
            I => \delay_measurement_inst.delay_tr_timer.N_287_4\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40780\,
            I => \delay_measurement_inst.delay_tr_timer.N_287_4\
        );

    \I__8839\ : InMux
    port map (
            O => \N__40775\,
            I => \N__40772\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__40772\,
            I => \N__40768\
        );

    \I__8837\ : InMux
    port map (
            O => \N__40771\,
            I => \N__40765\
        );

    \I__8836\ : Span4Mux_v
    port map (
            O => \N__40768\,
            I => \N__40761\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__40765\,
            I => \N__40758\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40764\,
            I => \N__40755\
        );

    \I__8833\ : Odrv4
    port map (
            O => \N__40761\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__8832\ : Odrv12
    port map (
            O => \N__40758\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__40755\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40748\,
            I => \N__40745\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__40745\,
            I => \N__40742\
        );

    \I__8828\ : Span4Mux_v
    port map (
            O => \N__40742\,
            I => \N__40738\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40735\
        );

    \I__8826\ : Odrv4
    port map (
            O => \N__40738\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__40735\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__8824\ : InMux
    port map (
            O => \N__40730\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__8823\ : CascadeMux
    port map (
            O => \N__40727\,
            I => \N__40724\
        );

    \I__8822\ : InMux
    port map (
            O => \N__40724\,
            I => \N__40721\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40721\,
            I => \N__40718\
        );

    \I__8820\ : Span4Mux_h
    port map (
            O => \N__40718\,
            I => \N__40714\
        );

    \I__8819\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40711\
        );

    \I__8818\ : Odrv4
    port map (
            O => \N__40714\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__40711\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40706\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__8815\ : CascadeMux
    port map (
            O => \N__40703\,
            I => \N__40697\
        );

    \I__8814\ : CascadeMux
    port map (
            O => \N__40702\,
            I => \N__40693\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40701\,
            I => \N__40687\
        );

    \I__8812\ : InMux
    port map (
            O => \N__40700\,
            I => \N__40680\
        );

    \I__8811\ : InMux
    port map (
            O => \N__40697\,
            I => \N__40680\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40696\,
            I => \N__40680\
        );

    \I__8809\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40675\
        );

    \I__8808\ : InMux
    port map (
            O => \N__40692\,
            I => \N__40675\
        );

    \I__8807\ : InMux
    port map (
            O => \N__40691\,
            I => \N__40672\
        );

    \I__8806\ : InMux
    port map (
            O => \N__40690\,
            I => \N__40669\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__40687\,
            I => \N__40666\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__40680\,
            I => \N__40661\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__40675\,
            I => \N__40661\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__40672\,
            I => \N__40656\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__40669\,
            I => \N__40656\
        );

    \I__8800\ : Span4Mux_h
    port map (
            O => \N__40666\,
            I => \N__40653\
        );

    \I__8799\ : Span4Mux_v
    port map (
            O => \N__40661\,
            I => \N__40650\
        );

    \I__8798\ : Span4Mux_h
    port map (
            O => \N__40656\,
            I => \N__40647\
        );

    \I__8797\ : Odrv4
    port map (
            O => \N__40653\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__8796\ : Odrv4
    port map (
            O => \N__40650\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__8795\ : Odrv4
    port map (
            O => \N__40647\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__8794\ : InMux
    port map (
            O => \N__40640\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__8793\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40634\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__40634\,
            I => \N__40631\
        );

    \I__8791\ : Span4Mux_v
    port map (
            O => \N__40631\,
            I => \N__40627\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40630\,
            I => \N__40624\
        );

    \I__8789\ : Span4Mux_v
    port map (
            O => \N__40627\,
            I => \N__40621\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__40624\,
            I => \N__40618\
        );

    \I__8787\ : Odrv4
    port map (
            O => \N__40621\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__8786\ : Odrv12
    port map (
            O => \N__40618\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40613\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__8784\ : CascadeMux
    port map (
            O => \N__40610\,
            I => \N__40606\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__40609\,
            I => \N__40603\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40598\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40603\,
            I => \N__40598\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__40598\,
            I => \N__40594\
        );

    \I__8779\ : InMux
    port map (
            O => \N__40597\,
            I => \N__40591\
        );

    \I__8778\ : Span4Mux_v
    port map (
            O => \N__40594\,
            I => \N__40588\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__40591\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__8776\ : Odrv4
    port map (
            O => \N__40588\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40583\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__8774\ : CascadeMux
    port map (
            O => \N__40580\,
            I => \N__40576\
        );

    \I__8773\ : CascadeMux
    port map (
            O => \N__40579\,
            I => \N__40573\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40567\
        );

    \I__8771\ : InMux
    port map (
            O => \N__40573\,
            I => \N__40567\
        );

    \I__8770\ : InMux
    port map (
            O => \N__40572\,
            I => \N__40564\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__40567\,
            I => \N__40561\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__40564\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__8767\ : Odrv12
    port map (
            O => \N__40561\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40556\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40553\,
            I => \N__40549\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40546\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__40549\,
            I => \N__40540\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__40546\,
            I => \N__40540\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40545\,
            I => \N__40537\
        );

    \I__8760\ : Span4Mux_v
    port map (
            O => \N__40540\,
            I => \N__40534\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__40537\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__8758\ : Odrv4
    port map (
            O => \N__40534\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__8757\ : InMux
    port map (
            O => \N__40529\,
            I => \bfn_15_28_0_\
        );

    \I__8756\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40522\
        );

    \I__8755\ : InMux
    port map (
            O => \N__40525\,
            I => \N__40519\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__40522\,
            I => \N__40513\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__40519\,
            I => \N__40513\
        );

    \I__8752\ : InMux
    port map (
            O => \N__40518\,
            I => \N__40510\
        );

    \I__8751\ : Span4Mux_v
    port map (
            O => \N__40513\,
            I => \N__40507\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__40510\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__8749\ : Odrv4
    port map (
            O => \N__40507\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40502\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__8747\ : CascadeMux
    port map (
            O => \N__40499\,
            I => \N__40495\
        );

    \I__8746\ : CascadeMux
    port map (
            O => \N__40498\,
            I => \N__40492\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40495\,
            I => \N__40487\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40492\,
            I => \N__40487\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__40487\,
            I => \N__40483\
        );

    \I__8742\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40480\
        );

    \I__8741\ : Span4Mux_h
    port map (
            O => \N__40483\,
            I => \N__40477\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__40480\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__8739\ : Odrv4
    port map (
            O => \N__40477\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__8738\ : InMux
    port map (
            O => \N__40472\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__8737\ : CascadeMux
    port map (
            O => \N__40469\,
            I => \N__40465\
        );

    \I__8736\ : CascadeMux
    port map (
            O => \N__40468\,
            I => \N__40462\
        );

    \I__8735\ : InMux
    port map (
            O => \N__40465\,
            I => \N__40457\
        );

    \I__8734\ : InMux
    port map (
            O => \N__40462\,
            I => \N__40457\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__40457\,
            I => \N__40453\
        );

    \I__8732\ : InMux
    port map (
            O => \N__40456\,
            I => \N__40450\
        );

    \I__8731\ : Span4Mux_h
    port map (
            O => \N__40453\,
            I => \N__40447\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__40450\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__8729\ : Odrv4
    port map (
            O => \N__40447\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__8728\ : InMux
    port map (
            O => \N__40442\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__8727\ : InMux
    port map (
            O => \N__40439\,
            I => \N__40436\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__40436\,
            I => \N__40432\
        );

    \I__8725\ : InMux
    port map (
            O => \N__40435\,
            I => \N__40429\
        );

    \I__8724\ : Span4Mux_h
    port map (
            O => \N__40432\,
            I => \N__40426\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__40429\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__8722\ : Odrv4
    port map (
            O => \N__40426\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__8721\ : InMux
    port map (
            O => \N__40421\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__8720\ : InMux
    port map (
            O => \N__40418\,
            I => \N__40396\
        );

    \I__8719\ : InMux
    port map (
            O => \N__40417\,
            I => \N__40396\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40416\,
            I => \N__40387\
        );

    \I__8717\ : InMux
    port map (
            O => \N__40415\,
            I => \N__40387\
        );

    \I__8716\ : InMux
    port map (
            O => \N__40414\,
            I => \N__40387\
        );

    \I__8715\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40387\
        );

    \I__8714\ : InMux
    port map (
            O => \N__40412\,
            I => \N__40366\
        );

    \I__8713\ : InMux
    port map (
            O => \N__40411\,
            I => \N__40366\
        );

    \I__8712\ : InMux
    port map (
            O => \N__40410\,
            I => \N__40366\
        );

    \I__8711\ : InMux
    port map (
            O => \N__40409\,
            I => \N__40366\
        );

    \I__8710\ : InMux
    port map (
            O => \N__40408\,
            I => \N__40357\
        );

    \I__8709\ : InMux
    port map (
            O => \N__40407\,
            I => \N__40357\
        );

    \I__8708\ : InMux
    port map (
            O => \N__40406\,
            I => \N__40357\
        );

    \I__8707\ : InMux
    port map (
            O => \N__40405\,
            I => \N__40357\
        );

    \I__8706\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40348\
        );

    \I__8705\ : InMux
    port map (
            O => \N__40403\,
            I => \N__40348\
        );

    \I__8704\ : InMux
    port map (
            O => \N__40402\,
            I => \N__40348\
        );

    \I__8703\ : InMux
    port map (
            O => \N__40401\,
            I => \N__40348\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__40396\,
            I => \N__40343\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__40387\,
            I => \N__40343\
        );

    \I__8700\ : InMux
    port map (
            O => \N__40386\,
            I => \N__40334\
        );

    \I__8699\ : InMux
    port map (
            O => \N__40385\,
            I => \N__40334\
        );

    \I__8698\ : InMux
    port map (
            O => \N__40384\,
            I => \N__40334\
        );

    \I__8697\ : InMux
    port map (
            O => \N__40383\,
            I => \N__40334\
        );

    \I__8696\ : InMux
    port map (
            O => \N__40382\,
            I => \N__40325\
        );

    \I__8695\ : InMux
    port map (
            O => \N__40381\,
            I => \N__40325\
        );

    \I__8694\ : InMux
    port map (
            O => \N__40380\,
            I => \N__40325\
        );

    \I__8693\ : InMux
    port map (
            O => \N__40379\,
            I => \N__40325\
        );

    \I__8692\ : InMux
    port map (
            O => \N__40378\,
            I => \N__40316\
        );

    \I__8691\ : InMux
    port map (
            O => \N__40377\,
            I => \N__40316\
        );

    \I__8690\ : InMux
    port map (
            O => \N__40376\,
            I => \N__40316\
        );

    \I__8689\ : InMux
    port map (
            O => \N__40375\,
            I => \N__40316\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__40366\,
            I => \N__40307\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__40357\,
            I => \N__40307\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__40348\,
            I => \N__40307\
        );

    \I__8685\ : Span4Mux_s3_v
    port map (
            O => \N__40343\,
            I => \N__40307\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__40334\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__40325\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__40316\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__40307\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__8680\ : InMux
    port map (
            O => \N__40298\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__8679\ : InMux
    port map (
            O => \N__40295\,
            I => \N__40292\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__40292\,
            I => \N__40288\
        );

    \I__8677\ : InMux
    port map (
            O => \N__40291\,
            I => \N__40285\
        );

    \I__8676\ : Span4Mux_h
    port map (
            O => \N__40288\,
            I => \N__40282\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__40285\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__8674\ : Odrv4
    port map (
            O => \N__40282\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__8673\ : CEMux
    port map (
            O => \N__40277\,
            I => \N__40265\
        );

    \I__8672\ : CEMux
    port map (
            O => \N__40276\,
            I => \N__40265\
        );

    \I__8671\ : CEMux
    port map (
            O => \N__40275\,
            I => \N__40265\
        );

    \I__8670\ : CEMux
    port map (
            O => \N__40274\,
            I => \N__40265\
        );

    \I__8669\ : GlobalMux
    port map (
            O => \N__40265\,
            I => \N__40262\
        );

    \I__8668\ : gio2CtrlBuf
    port map (
            O => \N__40262\,
            I => \current_shift_inst.timer_s1.N_181_i_g\
        );

    \I__8667\ : CascadeMux
    port map (
            O => \N__40259\,
            I => \N__40255\
        );

    \I__8666\ : CascadeMux
    port map (
            O => \N__40258\,
            I => \N__40252\
        );

    \I__8665\ : InMux
    port map (
            O => \N__40255\,
            I => \N__40246\
        );

    \I__8664\ : InMux
    port map (
            O => \N__40252\,
            I => \N__40246\
        );

    \I__8663\ : InMux
    port map (
            O => \N__40251\,
            I => \N__40243\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__40246\,
            I => \N__40240\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__40243\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__8660\ : Odrv12
    port map (
            O => \N__40240\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__8659\ : InMux
    port map (
            O => \N__40235\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__8658\ : CascadeMux
    port map (
            O => \N__40232\,
            I => \N__40228\
        );

    \I__8657\ : CascadeMux
    port map (
            O => \N__40231\,
            I => \N__40225\
        );

    \I__8656\ : InMux
    port map (
            O => \N__40228\,
            I => \N__40220\
        );

    \I__8655\ : InMux
    port map (
            O => \N__40225\,
            I => \N__40220\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__40220\,
            I => \N__40216\
        );

    \I__8653\ : InMux
    port map (
            O => \N__40219\,
            I => \N__40213\
        );

    \I__8652\ : Span4Mux_v
    port map (
            O => \N__40216\,
            I => \N__40210\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__40213\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__8650\ : Odrv4
    port map (
            O => \N__40210\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__8649\ : InMux
    port map (
            O => \N__40205\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__8648\ : InMux
    port map (
            O => \N__40202\,
            I => \N__40198\
        );

    \I__8647\ : InMux
    port map (
            O => \N__40201\,
            I => \N__40195\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__40198\,
            I => \N__40189\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__40195\,
            I => \N__40189\
        );

    \I__8644\ : InMux
    port map (
            O => \N__40194\,
            I => \N__40186\
        );

    \I__8643\ : Span4Mux_v
    port map (
            O => \N__40189\,
            I => \N__40183\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__40186\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__8641\ : Odrv4
    port map (
            O => \N__40183\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__8640\ : InMux
    port map (
            O => \N__40178\,
            I => \bfn_15_27_0_\
        );

    \I__8639\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40171\
        );

    \I__8638\ : InMux
    port map (
            O => \N__40174\,
            I => \N__40168\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__40171\,
            I => \N__40164\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__40168\,
            I => \N__40161\
        );

    \I__8635\ : InMux
    port map (
            O => \N__40167\,
            I => \N__40158\
        );

    \I__8634\ : Span4Mux_v
    port map (
            O => \N__40164\,
            I => \N__40153\
        );

    \I__8633\ : Span4Mux_v
    port map (
            O => \N__40161\,
            I => \N__40153\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__40158\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__8631\ : Odrv4
    port map (
            O => \N__40153\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__8630\ : InMux
    port map (
            O => \N__40148\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__8629\ : CascadeMux
    port map (
            O => \N__40145\,
            I => \N__40141\
        );

    \I__8628\ : CascadeMux
    port map (
            O => \N__40144\,
            I => \N__40138\
        );

    \I__8627\ : InMux
    port map (
            O => \N__40141\,
            I => \N__40133\
        );

    \I__8626\ : InMux
    port map (
            O => \N__40138\,
            I => \N__40133\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__40133\,
            I => \N__40129\
        );

    \I__8624\ : InMux
    port map (
            O => \N__40132\,
            I => \N__40126\
        );

    \I__8623\ : Span4Mux_h
    port map (
            O => \N__40129\,
            I => \N__40123\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__40126\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__8621\ : Odrv4
    port map (
            O => \N__40123\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__8620\ : InMux
    port map (
            O => \N__40118\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__8619\ : CascadeMux
    port map (
            O => \N__40115\,
            I => \N__40111\
        );

    \I__8618\ : CascadeMux
    port map (
            O => \N__40114\,
            I => \N__40108\
        );

    \I__8617\ : InMux
    port map (
            O => \N__40111\,
            I => \N__40103\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40108\,
            I => \N__40103\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__40103\,
            I => \N__40099\
        );

    \I__8614\ : InMux
    port map (
            O => \N__40102\,
            I => \N__40096\
        );

    \I__8613\ : Span4Mux_h
    port map (
            O => \N__40099\,
            I => \N__40093\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__40096\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__40093\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__8610\ : InMux
    port map (
            O => \N__40088\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40085\,
            I => \N__40078\
        );

    \I__8608\ : InMux
    port map (
            O => \N__40084\,
            I => \N__40078\
        );

    \I__8607\ : InMux
    port map (
            O => \N__40083\,
            I => \N__40075\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__40078\,
            I => \N__40072\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__40075\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__8604\ : Odrv12
    port map (
            O => \N__40072\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__8603\ : InMux
    port map (
            O => \N__40067\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__8602\ : InMux
    port map (
            O => \N__40064\,
            I => \N__40058\
        );

    \I__8601\ : InMux
    port map (
            O => \N__40063\,
            I => \N__40058\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__40058\,
            I => \N__40054\
        );

    \I__8599\ : InMux
    port map (
            O => \N__40057\,
            I => \N__40051\
        );

    \I__8598\ : Span4Mux_h
    port map (
            O => \N__40054\,
            I => \N__40048\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__40051\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__8596\ : Odrv4
    port map (
            O => \N__40048\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__8595\ : InMux
    port map (
            O => \N__40043\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__8594\ : InMux
    port map (
            O => \N__40040\,
            I => \N__40034\
        );

    \I__8593\ : InMux
    port map (
            O => \N__40039\,
            I => \N__40034\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__40034\,
            I => \N__40030\
        );

    \I__8591\ : InMux
    port map (
            O => \N__40033\,
            I => \N__40027\
        );

    \I__8590\ : Span4Mux_v
    port map (
            O => \N__40030\,
            I => \N__40024\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__40027\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__8588\ : Odrv4
    port map (
            O => \N__40024\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__8587\ : InMux
    port map (
            O => \N__40019\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__8586\ : InMux
    port map (
            O => \N__40016\,
            I => \N__40010\
        );

    \I__8585\ : InMux
    port map (
            O => \N__40015\,
            I => \N__40010\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__40010\,
            I => \N__40006\
        );

    \I__8583\ : InMux
    port map (
            O => \N__40009\,
            I => \N__40003\
        );

    \I__8582\ : Span4Mux_v
    port map (
            O => \N__40006\,
            I => \N__40000\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40003\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__8580\ : Odrv4
    port map (
            O => \N__40000\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__8579\ : InMux
    port map (
            O => \N__39995\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__8578\ : CascadeMux
    port map (
            O => \N__39992\,
            I => \N__39988\
        );

    \I__8577\ : InMux
    port map (
            O => \N__39991\,
            I => \N__39985\
        );

    \I__8576\ : InMux
    port map (
            O => \N__39988\,
            I => \N__39982\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__39985\,
            I => \N__39976\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__39982\,
            I => \N__39976\
        );

    \I__8573\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39973\
        );

    \I__8572\ : Span4Mux_v
    port map (
            O => \N__39976\,
            I => \N__39970\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__39973\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__8570\ : Odrv4
    port map (
            O => \N__39970\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__8569\ : InMux
    port map (
            O => \N__39965\,
            I => \bfn_15_26_0_\
        );

    \I__8568\ : CascadeMux
    port map (
            O => \N__39962\,
            I => \N__39958\
        );

    \I__8567\ : InMux
    port map (
            O => \N__39961\,
            I => \N__39955\
        );

    \I__8566\ : InMux
    port map (
            O => \N__39958\,
            I => \N__39952\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__39955\,
            I => \N__39946\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__39952\,
            I => \N__39946\
        );

    \I__8563\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39943\
        );

    \I__8562\ : Span4Mux_v
    port map (
            O => \N__39946\,
            I => \N__39940\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__39943\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__8560\ : Odrv4
    port map (
            O => \N__39940\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__8559\ : InMux
    port map (
            O => \N__39935\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__8558\ : CascadeMux
    port map (
            O => \N__39932\,
            I => \N__39928\
        );

    \I__8557\ : CascadeMux
    port map (
            O => \N__39931\,
            I => \N__39925\
        );

    \I__8556\ : InMux
    port map (
            O => \N__39928\,
            I => \N__39920\
        );

    \I__8555\ : InMux
    port map (
            O => \N__39925\,
            I => \N__39920\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__39920\,
            I => \N__39916\
        );

    \I__8553\ : InMux
    port map (
            O => \N__39919\,
            I => \N__39913\
        );

    \I__8552\ : Span4Mux_h
    port map (
            O => \N__39916\,
            I => \N__39910\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__39913\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__8550\ : Odrv4
    port map (
            O => \N__39910\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__8549\ : InMux
    port map (
            O => \N__39905\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__8548\ : CascadeMux
    port map (
            O => \N__39902\,
            I => \N__39898\
        );

    \I__8547\ : CascadeMux
    port map (
            O => \N__39901\,
            I => \N__39895\
        );

    \I__8546\ : InMux
    port map (
            O => \N__39898\,
            I => \N__39889\
        );

    \I__8545\ : InMux
    port map (
            O => \N__39895\,
            I => \N__39889\
        );

    \I__8544\ : InMux
    port map (
            O => \N__39894\,
            I => \N__39886\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__39889\,
            I => \N__39883\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__39886\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__8541\ : Odrv12
    port map (
            O => \N__39883\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__8540\ : InMux
    port map (
            O => \N__39878\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__8539\ : InMux
    port map (
            O => \N__39875\,
            I => \N__39868\
        );

    \I__8538\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39868\
        );

    \I__8537\ : InMux
    port map (
            O => \N__39873\,
            I => \N__39865\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__39868\,
            I => \N__39862\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__39865\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__8534\ : Odrv12
    port map (
            O => \N__39862\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__8533\ : InMux
    port map (
            O => \N__39857\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__8532\ : InMux
    port map (
            O => \N__39854\,
            I => \N__39847\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39853\,
            I => \N__39847\
        );

    \I__8530\ : InMux
    port map (
            O => \N__39852\,
            I => \N__39844\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__39847\,
            I => \N__39841\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__39844\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__8527\ : Odrv12
    port map (
            O => \N__39841\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__8526\ : InMux
    port map (
            O => \N__39836\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39833\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39830\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__8523\ : InMux
    port map (
            O => \N__39827\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__8522\ : InMux
    port map (
            O => \N__39824\,
            I => \bfn_15_25_0_\
        );

    \I__8521\ : InMux
    port map (
            O => \N__39821\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__8520\ : InMux
    port map (
            O => \N__39818\,
            I => \N__39811\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39817\,
            I => \N__39811\
        );

    \I__8518\ : InMux
    port map (
            O => \N__39816\,
            I => \N__39808\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__39811\,
            I => \N__39805\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__39808\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__8515\ : Odrv12
    port map (
            O => \N__39805\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__8514\ : InMux
    port map (
            O => \N__39800\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__8513\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39791\
        );

    \I__8512\ : InMux
    port map (
            O => \N__39796\,
            I => \N__39791\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__39791\,
            I => \N__39787\
        );

    \I__8510\ : InMux
    port map (
            O => \N__39790\,
            I => \N__39784\
        );

    \I__8509\ : Span4Mux_h
    port map (
            O => \N__39787\,
            I => \N__39781\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__39784\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__8507\ : Odrv4
    port map (
            O => \N__39781\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39776\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__8505\ : CascadeMux
    port map (
            O => \N__39773\,
            I => \N__39769\
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__39772\,
            I => \N__39766\
        );

    \I__8503\ : InMux
    port map (
            O => \N__39769\,
            I => \N__39760\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39766\,
            I => \N__39760\
        );

    \I__8501\ : InMux
    port map (
            O => \N__39765\,
            I => \N__39757\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__39760\,
            I => \N__39754\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__39757\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__8498\ : Odrv12
    port map (
            O => \N__39754\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__8497\ : InMux
    port map (
            O => \N__39749\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__8496\ : CascadeMux
    port map (
            O => \N__39746\,
            I => \N__39742\
        );

    \I__8495\ : CascadeMux
    port map (
            O => \N__39745\,
            I => \N__39739\
        );

    \I__8494\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39733\
        );

    \I__8493\ : InMux
    port map (
            O => \N__39739\,
            I => \N__39733\
        );

    \I__8492\ : InMux
    port map (
            O => \N__39738\,
            I => \N__39730\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__39733\,
            I => \N__39727\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__39730\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__8489\ : Odrv12
    port map (
            O => \N__39727\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__8488\ : InMux
    port map (
            O => \N__39722\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39719\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__8486\ : InMux
    port map (
            O => \N__39716\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__8485\ : InMux
    port map (
            O => \N__39713\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__8484\ : InMux
    port map (
            O => \N__39710\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__8483\ : InMux
    port map (
            O => \N__39707\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__8482\ : InMux
    port map (
            O => \N__39704\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39701\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__8480\ : InMux
    port map (
            O => \N__39698\,
            I => \bfn_15_24_0_\
        );

    \I__8479\ : InMux
    port map (
            O => \N__39695\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__8478\ : InMux
    port map (
            O => \N__39692\,
            I => \bfn_15_22_0_\
        );

    \I__8477\ : InMux
    port map (
            O => \N__39689\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__8476\ : InMux
    port map (
            O => \N__39686\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__8475\ : InMux
    port map (
            O => \N__39683\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__8474\ : InMux
    port map (
            O => \N__39680\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__8473\ : InMux
    port map (
            O => \N__39677\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__8472\ : InMux
    port map (
            O => \N__39674\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39671\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39668\,
            I => \bfn_15_23_0_\
        );

    \I__8469\ : InMux
    port map (
            O => \N__39665\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__8468\ : InMux
    port map (
            O => \N__39662\,
            I => \N__39659\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__39659\,
            I => \N__39656\
        );

    \I__8466\ : Span4Mux_h
    port map (
            O => \N__39656\,
            I => \N__39653\
        );

    \I__8465\ : Odrv4
    port map (
            O => \N__39653\,
            I => \current_shift_inst.control_input_1_axb_11\
        );

    \I__8464\ : InMux
    port map (
            O => \N__39650\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__8463\ : InMux
    port map (
            O => \N__39647\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__8462\ : InMux
    port map (
            O => \N__39644\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__8461\ : InMux
    port map (
            O => \N__39641\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39638\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39635\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__8458\ : InMux
    port map (
            O => \N__39632\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__8457\ : CascadeMux
    port map (
            O => \N__39629\,
            I => \N__39626\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39626\,
            I => \N__39623\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__39623\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__8454\ : InMux
    port map (
            O => \N__39620\,
            I => \N__39617\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__39617\,
            I => \N__39614\
        );

    \I__8452\ : Span4Mux_v
    port map (
            O => \N__39614\,
            I => \N__39611\
        );

    \I__8451\ : Odrv4
    port map (
            O => \N__39611\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39608\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39605\,
            I => \N__39602\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39602\,
            I => \N__39599\
        );

    \I__8447\ : Span4Mux_h
    port map (
            O => \N__39599\,
            I => \N__39596\
        );

    \I__8446\ : Odrv4
    port map (
            O => \N__39596\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__8445\ : InMux
    port map (
            O => \N__39593\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__8444\ : CascadeMux
    port map (
            O => \N__39590\,
            I => \N__39587\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39587\,
            I => \N__39584\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__39584\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39581\,
            I => \N__39578\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__39578\,
            I => \N__39575\
        );

    \I__8439\ : Span4Mux_h
    port map (
            O => \N__39575\,
            I => \N__39572\
        );

    \I__8438\ : Odrv4
    port map (
            O => \N__39572\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__8437\ : InMux
    port map (
            O => \N__39569\,
            I => \bfn_15_20_0_\
        );

    \I__8436\ : InMux
    port map (
            O => \N__39566\,
            I => \N__39563\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__39563\,
            I => \N__39560\
        );

    \I__8434\ : Span4Mux_h
    port map (
            O => \N__39560\,
            I => \N__39557\
        );

    \I__8433\ : Odrv4
    port map (
            O => \N__39557\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__8432\ : InMux
    port map (
            O => \N__39554\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__8431\ : InMux
    port map (
            O => \N__39551\,
            I => \N__39548\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__39548\,
            I => \N__39545\
        );

    \I__8429\ : Span4Mux_h
    port map (
            O => \N__39545\,
            I => \N__39542\
        );

    \I__8428\ : Odrv4
    port map (
            O => \N__39542\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39539\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39536\,
            I => \N__39533\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__39533\,
            I => \N__39530\
        );

    \I__8424\ : Span4Mux_v
    port map (
            O => \N__39530\,
            I => \N__39527\
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__39527\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__8422\ : InMux
    port map (
            O => \N__39524\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__8421\ : InMux
    port map (
            O => \N__39521\,
            I => \N__39518\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__39518\,
            I => \N__39515\
        );

    \I__8419\ : Odrv4
    port map (
            O => \N__39515\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__8418\ : InMux
    port map (
            O => \N__39512\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__8417\ : InMux
    port map (
            O => \N__39509\,
            I => \N__39506\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__39506\,
            I => \N__39503\
        );

    \I__8415\ : Odrv12
    port map (
            O => \N__39503\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__8414\ : InMux
    port map (
            O => \N__39500\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39497\,
            I => \N__39494\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__39494\,
            I => \N__39491\
        );

    \I__8411\ : Odrv12
    port map (
            O => \N__39491\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__8410\ : InMux
    port map (
            O => \N__39488\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39485\,
            I => \N__39482\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__39482\,
            I => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\
        );

    \I__8407\ : InMux
    port map (
            O => \N__39479\,
            I => \N__39476\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__39476\,
            I => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__39473\,
            I => \N__39470\
        );

    \I__8404\ : InMux
    port map (
            O => \N__39470\,
            I => \N__39467\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__39467\,
            I => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\
        );

    \I__8402\ : InMux
    port map (
            O => \N__39464\,
            I => \N__39461\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__39461\,
            I => \N__39458\
        );

    \I__8400\ : Odrv4
    port map (
            O => \N__39458\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__8399\ : InMux
    port map (
            O => \N__39455\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__8398\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39449\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__39449\,
            I => \N__39446\
        );

    \I__8396\ : Odrv12
    port map (
            O => \N__39446\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__8395\ : InMux
    port map (
            O => \N__39443\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__8394\ : InMux
    port map (
            O => \N__39440\,
            I => \N__39437\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__39437\,
            I => \N__39434\
        );

    \I__8392\ : Span4Mux_v
    port map (
            O => \N__39434\,
            I => \N__39431\
        );

    \I__8391\ : Odrv4
    port map (
            O => \N__39431\,
            I => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\
        );

    \I__8390\ : InMux
    port map (
            O => \N__39428\,
            I => \N__39425\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__39425\,
            I => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\
        );

    \I__8388\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39419\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__39419\,
            I => \N__39416\
        );

    \I__8386\ : Odrv12
    port map (
            O => \N__39416\,
            I => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\
        );

    \I__8385\ : InMux
    port map (
            O => \N__39413\,
            I => \N__39410\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__39410\,
            I => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\
        );

    \I__8383\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39404\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__39404\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__8381\ : InMux
    port map (
            O => \N__39401\,
            I => \N__39398\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__39398\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__8379\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39392\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__39392\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__8377\ : InMux
    port map (
            O => \N__39389\,
            I => \N__39386\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__39386\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__8375\ : InMux
    port map (
            O => \N__39383\,
            I => \N__39380\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__39380\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39374\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__39374\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__8371\ : CascadeMux
    port map (
            O => \N__39371\,
            I => \N__39368\
        );

    \I__8370\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39365\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__39365\,
            I => \N__39362\
        );

    \I__8368\ : Odrv4
    port map (
            O => \N__39362\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39359\,
            I => \N__39356\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__39356\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__8365\ : InMux
    port map (
            O => \N__39353\,
            I => \N__39350\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__39350\,
            I => \N__39347\
        );

    \I__8363\ : Odrv4
    port map (
            O => \N__39347\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__8362\ : CascadeMux
    port map (
            O => \N__39344\,
            I => \N__39341\
        );

    \I__8361\ : InMux
    port map (
            O => \N__39341\,
            I => \N__39338\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__39338\,
            I => \N__39335\
        );

    \I__8359\ : Odrv4
    port map (
            O => \N__39335\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__8358\ : InMux
    port map (
            O => \N__39332\,
            I => \N__39328\
        );

    \I__8357\ : InMux
    port map (
            O => \N__39331\,
            I => \N__39323\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__39328\,
            I => \N__39320\
        );

    \I__8355\ : InMux
    port map (
            O => \N__39327\,
            I => \N__39317\
        );

    \I__8354\ : CascadeMux
    port map (
            O => \N__39326\,
            I => \N__39314\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__39323\,
            I => \N__39311\
        );

    \I__8352\ : Span4Mux_h
    port map (
            O => \N__39320\,
            I => \N__39308\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__39317\,
            I => \N__39305\
        );

    \I__8350\ : InMux
    port map (
            O => \N__39314\,
            I => \N__39302\
        );

    \I__8349\ : Span4Mux_v
    port map (
            O => \N__39311\,
            I => \N__39297\
        );

    \I__8348\ : Span4Mux_v
    port map (
            O => \N__39308\,
            I => \N__39297\
        );

    \I__8347\ : Span12Mux_v
    port map (
            O => \N__39305\,
            I => \N__39294\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__39302\,
            I => measured_delay_tr_7
        );

    \I__8345\ : Odrv4
    port map (
            O => \N__39297\,
            I => measured_delay_tr_7
        );

    \I__8344\ : Odrv12
    port map (
            O => \N__39294\,
            I => measured_delay_tr_7
        );

    \I__8343\ : InMux
    port map (
            O => \N__39287\,
            I => \N__39281\
        );

    \I__8342\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39281\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__39281\,
            I => \N__39278\
        );

    \I__8340\ : Span4Mux_v
    port map (
            O => \N__39278\,
            I => \N__39274\
        );

    \I__8339\ : InMux
    port map (
            O => \N__39277\,
            I => \N__39271\
        );

    \I__8338\ : Span4Mux_v
    port map (
            O => \N__39274\,
            I => \N__39268\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__39271\,
            I => \N__39265\
        );

    \I__8336\ : Odrv4
    port map (
            O => \N__39268\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i\
        );

    \I__8335\ : Odrv4
    port map (
            O => \N__39265\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i\
        );

    \I__8334\ : CascadeMux
    port map (
            O => \N__39260\,
            I => \N__39256\
        );

    \I__8333\ : CascadeMux
    port map (
            O => \N__39259\,
            I => \N__39253\
        );

    \I__8332\ : InMux
    port map (
            O => \N__39256\,
            I => \N__39244\
        );

    \I__8331\ : InMux
    port map (
            O => \N__39253\,
            I => \N__39237\
        );

    \I__8330\ : InMux
    port map (
            O => \N__39252\,
            I => \N__39237\
        );

    \I__8329\ : InMux
    port map (
            O => \N__39251\,
            I => \N__39237\
        );

    \I__8328\ : InMux
    port map (
            O => \N__39250\,
            I => \N__39232\
        );

    \I__8327\ : InMux
    port map (
            O => \N__39249\,
            I => \N__39232\
        );

    \I__8326\ : InMux
    port map (
            O => \N__39248\,
            I => \N__39227\
        );

    \I__8325\ : InMux
    port map (
            O => \N__39247\,
            I => \N__39227\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__39244\,
            I => \N__39220\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__39237\,
            I => \N__39220\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39232\,
            I => \N__39220\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__39227\,
            I => \N__39217\
        );

    \I__8320\ : Span4Mux_v
    port map (
            O => \N__39220\,
            I => \N__39214\
        );

    \I__8319\ : Span12Mux_v
    port map (
            O => \N__39217\,
            I => \N__39211\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__39214\,
            I => \delay_measurement_inst.N_267\
        );

    \I__8317\ : Odrv12
    port map (
            O => \N__39211\,
            I => \delay_measurement_inst.N_267\
        );

    \I__8316\ : InMux
    port map (
            O => \N__39206\,
            I => \N__39201\
        );

    \I__8315\ : InMux
    port map (
            O => \N__39205\,
            I => \N__39198\
        );

    \I__8314\ : InMux
    port map (
            O => \N__39204\,
            I => \N__39195\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__39201\,
            I => \N__39190\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__39198\,
            I => \N__39190\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__39195\,
            I => \N__39184\
        );

    \I__8310\ : Span4Mux_h
    port map (
            O => \N__39190\,
            I => \N__39184\
        );

    \I__8309\ : CascadeMux
    port map (
            O => \N__39189\,
            I => \N__39181\
        );

    \I__8308\ : Span4Mux_v
    port map (
            O => \N__39184\,
            I => \N__39178\
        );

    \I__8307\ : InMux
    port map (
            O => \N__39181\,
            I => \N__39175\
        );

    \I__8306\ : Span4Mux_v
    port map (
            O => \N__39178\,
            I => \N__39172\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__39175\,
            I => measured_delay_tr_8
        );

    \I__8304\ : Odrv4
    port map (
            O => \N__39172\,
            I => measured_delay_tr_8
        );

    \I__8303\ : InMux
    port map (
            O => \N__39167\,
            I => \N__39164\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__39164\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__8301\ : CascadeMux
    port map (
            O => \N__39161\,
            I => \N__39157\
        );

    \I__8300\ : InMux
    port map (
            O => \N__39160\,
            I => \N__39154\
        );

    \I__8299\ : InMux
    port map (
            O => \N__39157\,
            I => \N__39151\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__39154\,
            I => \current_shift_inst.N_1318_i\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__39151\,
            I => \current_shift_inst.N_1318_i\
        );

    \I__8296\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39143\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__39143\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__8294\ : InMux
    port map (
            O => \N__39140\,
            I => \N__39137\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__39137\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__8292\ : InMux
    port map (
            O => \N__39134\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__8291\ : InMux
    port map (
            O => \N__39131\,
            I => \N__39128\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__39128\,
            I => \N__39124\
        );

    \I__8289\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39121\
        );

    \I__8288\ : Span4Mux_v
    port map (
            O => \N__39124\,
            I => \N__39118\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__39121\,
            I => \N__39115\
        );

    \I__8286\ : Span4Mux_v
    port map (
            O => \N__39118\,
            I => \N__39110\
        );

    \I__8285\ : Span4Mux_v
    port map (
            O => \N__39115\,
            I => \N__39107\
        );

    \I__8284\ : InMux
    port map (
            O => \N__39114\,
            I => \N__39104\
        );

    \I__8283\ : InMux
    port map (
            O => \N__39113\,
            I => \N__39101\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__39110\,
            I => measured_delay_tr_17
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__39107\,
            I => measured_delay_tr_17
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__39104\,
            I => measured_delay_tr_17
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__39101\,
            I => measured_delay_tr_17
        );

    \I__8278\ : CascadeMux
    port map (
            O => \N__39092\,
            I => \N__39089\
        );

    \I__8277\ : InMux
    port map (
            O => \N__39089\,
            I => \N__39086\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__39086\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__8275\ : InMux
    port map (
            O => \N__39083\,
            I => \N__39080\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__39080\,
            I => \N__39076\
        );

    \I__8273\ : InMux
    port map (
            O => \N__39079\,
            I => \N__39073\
        );

    \I__8272\ : Span4Mux_v
    port map (
            O => \N__39076\,
            I => \N__39067\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__39073\,
            I => \N__39067\
        );

    \I__8270\ : InMux
    port map (
            O => \N__39072\,
            I => \N__39064\
        );

    \I__8269\ : Span4Mux_h
    port map (
            O => \N__39067\,
            I => \N__39060\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__39064\,
            I => \N__39057\
        );

    \I__8267\ : InMux
    port map (
            O => \N__39063\,
            I => \N__39054\
        );

    \I__8266\ : Odrv4
    port map (
            O => \N__39060\,
            I => measured_delay_tr_18
        );

    \I__8265\ : Odrv4
    port map (
            O => \N__39057\,
            I => measured_delay_tr_18
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__39054\,
            I => measured_delay_tr_18
        );

    \I__8263\ : CascadeMux
    port map (
            O => \N__39047\,
            I => \N__39044\
        );

    \I__8262\ : InMux
    port map (
            O => \N__39044\,
            I => \N__39041\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__39041\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__8260\ : CEMux
    port map (
            O => \N__39038\,
            I => \N__39033\
        );

    \I__8259\ : CEMux
    port map (
            O => \N__39037\,
            I => \N__39030\
        );

    \I__8258\ : CEMux
    port map (
            O => \N__39036\,
            I => \N__39027\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__39033\,
            I => \N__39023\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__39030\,
            I => \N__39020\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__39027\,
            I => \N__39017\
        );

    \I__8254\ : CEMux
    port map (
            O => \N__39026\,
            I => \N__39014\
        );

    \I__8253\ : Odrv4
    port map (
            O => \N__39023\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__39020\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__8251\ : Odrv12
    port map (
            O => \N__39017\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__39014\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__8249\ : CascadeMux
    port map (
            O => \N__39005\,
            I => \N__39002\
        );

    \I__8248\ : InMux
    port map (
            O => \N__39002\,
            I => \N__38999\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__38999\,
            I => \N__38996\
        );

    \I__8246\ : Odrv4
    port map (
            O => \N__38996\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__8245\ : InMux
    port map (
            O => \N__38993\,
            I => \N__38990\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__38990\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__8243\ : CascadeMux
    port map (
            O => \N__38987\,
            I => \N__38984\
        );

    \I__8242\ : InMux
    port map (
            O => \N__38984\,
            I => \N__38981\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__38981\,
            I => \N__38978\
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__38978\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__8239\ : InMux
    port map (
            O => \N__38975\,
            I => \N__38972\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__38972\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__8237\ : CascadeMux
    port map (
            O => \N__38969\,
            I => \N__38966\
        );

    \I__8236\ : InMux
    port map (
            O => \N__38966\,
            I => \N__38963\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__38963\,
            I => \N__38960\
        );

    \I__8234\ : Span4Mux_v
    port map (
            O => \N__38960\,
            I => \N__38957\
        );

    \I__8233\ : Odrv4
    port map (
            O => \N__38957\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__8232\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38951\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__38951\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__8230\ : CascadeMux
    port map (
            O => \N__38948\,
            I => \N__38945\
        );

    \I__8229\ : InMux
    port map (
            O => \N__38945\,
            I => \N__38942\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__38942\,
            I => \N__38939\
        );

    \I__8227\ : Odrv4
    port map (
            O => \N__38939\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__8226\ : InMux
    port map (
            O => \N__38936\,
            I => \N__38933\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__38933\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__8224\ : CascadeMux
    port map (
            O => \N__38930\,
            I => \N__38927\
        );

    \I__8223\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38924\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__38924\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__8221\ : InMux
    port map (
            O => \N__38921\,
            I => \N__38918\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__38918\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__8219\ : InMux
    port map (
            O => \N__38915\,
            I => \N__38912\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__38912\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__8217\ : InMux
    port map (
            O => \N__38909\,
            I => \N__38906\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__38906\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__8215\ : CascadeMux
    port map (
            O => \N__38903\,
            I => \N__38900\
        );

    \I__8214\ : InMux
    port map (
            O => \N__38900\,
            I => \N__38897\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__38897\,
            I => \N__38894\
        );

    \I__8212\ : Span4Mux_h
    port map (
            O => \N__38894\,
            I => \N__38891\
        );

    \I__8211\ : Odrv4
    port map (
            O => \N__38891\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__8210\ : InMux
    port map (
            O => \N__38888\,
            I => \N__38885\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__38885\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__38882\,
            I => \N__38879\
        );

    \I__8207\ : InMux
    port map (
            O => \N__38879\,
            I => \N__38876\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__38876\,
            I => \N__38873\
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__38873\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__8204\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38867\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__38867\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__8202\ : CascadeMux
    port map (
            O => \N__38864\,
            I => \N__38861\
        );

    \I__8201\ : InMux
    port map (
            O => \N__38861\,
            I => \N__38858\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__38858\,
            I => \N__38855\
        );

    \I__8199\ : Odrv4
    port map (
            O => \N__38855\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__8198\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38849\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__38849\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__8196\ : CascadeMux
    port map (
            O => \N__38846\,
            I => \N__38843\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38843\,
            I => \N__38840\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__38840\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__8193\ : InMux
    port map (
            O => \N__38837\,
            I => \N__38834\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__38834\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__8191\ : CascadeMux
    port map (
            O => \N__38831\,
            I => \N__38828\
        );

    \I__8190\ : InMux
    port map (
            O => \N__38828\,
            I => \N__38825\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__38825\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38819\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__38819\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__38816\,
            I => \N__38813\
        );

    \I__8185\ : InMux
    port map (
            O => \N__38813\,
            I => \N__38810\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__38810\,
            I => \N__38807\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__38807\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__8182\ : InMux
    port map (
            O => \N__38804\,
            I => \N__38801\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__38801\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__38798\,
            I => \N__38795\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38795\,
            I => \N__38792\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__38792\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__8177\ : InMux
    port map (
            O => \N__38789\,
            I => \N__38786\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38786\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__8175\ : CascadeMux
    port map (
            O => \N__38783\,
            I => \N__38780\
        );

    \I__8174\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38777\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__38777\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38771\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__38771\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__8170\ : CascadeMux
    port map (
            O => \N__38768\,
            I => \N__38765\
        );

    \I__8169\ : InMux
    port map (
            O => \N__38765\,
            I => \N__38762\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__38762\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__8167\ : InMux
    port map (
            O => \N__38759\,
            I => \N__38756\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__38756\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38753\,
            I => \N__38750\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__38750\,
            I => \N__38744\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38749\,
            I => \N__38741\
        );

    \I__8162\ : CascadeMux
    port map (
            O => \N__38748\,
            I => \N__38738\
        );

    \I__8161\ : CascadeMux
    port map (
            O => \N__38747\,
            I => \N__38735\
        );

    \I__8160\ : Span4Mux_v
    port map (
            O => \N__38744\,
            I => \N__38730\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38741\,
            I => \N__38730\
        );

    \I__8158\ : InMux
    port map (
            O => \N__38738\,
            I => \N__38727\
        );

    \I__8157\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38724\
        );

    \I__8156\ : Odrv4
    port map (
            O => \N__38730\,
            I => measured_delay_tr_19
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__38727\,
            I => measured_delay_tr_19
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38724\,
            I => measured_delay_tr_19
        );

    \I__8153\ : InMux
    port map (
            O => \N__38717\,
            I => \N__38714\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__38714\,
            I => \N__38710\
        );

    \I__8151\ : InMux
    port map (
            O => \N__38713\,
            I => \N__38707\
        );

    \I__8150\ : Span4Mux_h
    port map (
            O => \N__38710\,
            I => \N__38701\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__38707\,
            I => \N__38701\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38706\,
            I => \N__38698\
        );

    \I__8147\ : Odrv4
    port map (
            O => \N__38701\,
            I => measured_delay_tr_12
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__38698\,
            I => measured_delay_tr_12
        );

    \I__8145\ : InMux
    port map (
            O => \N__38693\,
            I => \N__38689\
        );

    \I__8144\ : InMux
    port map (
            O => \N__38692\,
            I => \N__38683\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__38689\,
            I => \N__38680\
        );

    \I__8142\ : InMux
    port map (
            O => \N__38688\,
            I => \N__38677\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38687\,
            I => \N__38672\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38686\,
            I => \N__38672\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__38683\,
            I => \N__38669\
        );

    \I__8138\ : Span4Mux_h
    port map (
            O => \N__38680\,
            I => \N__38664\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__38677\,
            I => \N__38664\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__38672\,
            I => \N__38661\
        );

    \I__8135\ : Span4Mux_h
    port map (
            O => \N__38669\,
            I => \N__38658\
        );

    \I__8134\ : Span4Mux_v
    port map (
            O => \N__38664\,
            I => \N__38655\
        );

    \I__8133\ : Span4Mux_h
    port map (
            O => \N__38661\,
            I => \N__38652\
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__38658\,
            I => measured_delay_tr_14
        );

    \I__8131\ : Odrv4
    port map (
            O => \N__38655\,
            I => measured_delay_tr_14
        );

    \I__8130\ : Odrv4
    port map (
            O => \N__38652\,
            I => measured_delay_tr_14
        );

    \I__8129\ : InMux
    port map (
            O => \N__38645\,
            I => \N__38636\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38644\,
            I => \N__38636\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38643\,
            I => \N__38631\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38642\,
            I => \N__38631\
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__38641\,
            I => \N__38628\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38636\,
            I => \N__38623\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__38631\,
            I => \N__38620\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38628\,
            I => \N__38613\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38627\,
            I => \N__38613\
        );

    \I__8120\ : InMux
    port map (
            O => \N__38626\,
            I => \N__38613\
        );

    \I__8119\ : Span4Mux_h
    port map (
            O => \N__38623\,
            I => \N__38608\
        );

    \I__8118\ : Span4Mux_h
    port map (
            O => \N__38620\,
            I => \N__38603\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__38613\,
            I => \N__38603\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38612\,
            I => \N__38598\
        );

    \I__8115\ : InMux
    port map (
            O => \N__38611\,
            I => \N__38598\
        );

    \I__8114\ : Odrv4
    port map (
            O => \N__38608\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__38603\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__38598\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__8111\ : InMux
    port map (
            O => \N__38591\,
            I => \N__38587\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38584\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__38587\,
            I => \N__38580\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__38584\,
            I => \N__38577\
        );

    \I__8107\ : CascadeMux
    port map (
            O => \N__38583\,
            I => \N__38574\
        );

    \I__8106\ : Span4Mux_v
    port map (
            O => \N__38580\,
            I => \N__38571\
        );

    \I__8105\ : Span4Mux_h
    port map (
            O => \N__38577\,
            I => \N__38568\
        );

    \I__8104\ : InMux
    port map (
            O => \N__38574\,
            I => \N__38565\
        );

    \I__8103\ : Odrv4
    port map (
            O => \N__38571\,
            I => measured_delay_tr_13
        );

    \I__8102\ : Odrv4
    port map (
            O => \N__38568\,
            I => measured_delay_tr_13
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__38565\,
            I => measured_delay_tr_13
        );

    \I__8100\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38552\
        );

    \I__8099\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38552\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__38552\,
            I => \N__38546\
        );

    \I__8097\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38542\
        );

    \I__8096\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38539\
        );

    \I__8095\ : InMux
    port map (
            O => \N__38549\,
            I => \N__38536\
        );

    \I__8094\ : Span4Mux_v
    port map (
            O => \N__38546\,
            I => \N__38533\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38545\,
            I => \N__38530\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__38542\,
            I => \N__38527\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__38539\,
            I => \N__38524\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__38536\,
            I => \N__38521\
        );

    \I__8089\ : Span4Mux_v
    port map (
            O => \N__38533\,
            I => \N__38516\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__38530\,
            I => \N__38516\
        );

    \I__8087\ : Span4Mux_v
    port map (
            O => \N__38527\,
            I => \N__38513\
        );

    \I__8086\ : Span4Mux_h
    port map (
            O => \N__38524\,
            I => \N__38506\
        );

    \I__8085\ : Span4Mux_v
    port map (
            O => \N__38521\,
            I => \N__38506\
        );

    \I__8084\ : Span4Mux_h
    port map (
            O => \N__38516\,
            I => \N__38506\
        );

    \I__8083\ : Odrv4
    port map (
            O => \N__38513\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__8082\ : Odrv4
    port map (
            O => \N__38506\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__8081\ : InMux
    port map (
            O => \N__38501\,
            I => \N__38492\
        );

    \I__8080\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38492\
        );

    \I__8079\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38489\
        );

    \I__8078\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38485\
        );

    \I__8077\ : InMux
    port map (
            O => \N__38497\,
            I => \N__38482\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__38492\,
            I => \N__38479\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__38489\,
            I => \N__38476\
        );

    \I__8074\ : InMux
    port map (
            O => \N__38488\,
            I => \N__38473\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__38485\,
            I => \N__38468\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__38482\,
            I => \N__38463\
        );

    \I__8071\ : Span4Mux_h
    port map (
            O => \N__38479\,
            I => \N__38463\
        );

    \I__8070\ : Span4Mux_h
    port map (
            O => \N__38476\,
            I => \N__38457\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__38473\,
            I => \N__38457\
        );

    \I__8068\ : InMux
    port map (
            O => \N__38472\,
            I => \N__38454\
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__38471\,
            I => \N__38450\
        );

    \I__8066\ : Span4Mux_v
    port map (
            O => \N__38468\,
            I => \N__38447\
        );

    \I__8065\ : Span4Mux_v
    port map (
            O => \N__38463\,
            I => \N__38444\
        );

    \I__8064\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38441\
        );

    \I__8063\ : Sp12to4
    port map (
            O => \N__38457\,
            I => \N__38436\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__38454\,
            I => \N__38436\
        );

    \I__8061\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38431\
        );

    \I__8060\ : InMux
    port map (
            O => \N__38450\,
            I => \N__38431\
        );

    \I__8059\ : Odrv4
    port map (
            O => \N__38447\,
            I => measured_delay_tr_15
        );

    \I__8058\ : Odrv4
    port map (
            O => \N__38444\,
            I => measured_delay_tr_15
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__38441\,
            I => measured_delay_tr_15
        );

    \I__8056\ : Odrv12
    port map (
            O => \N__38436\,
            I => measured_delay_tr_15
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__38431\,
            I => measured_delay_tr_15
        );

    \I__8054\ : CascadeMux
    port map (
            O => \N__38420\,
            I => \N__38417\
        );

    \I__8053\ : InMux
    port map (
            O => \N__38417\,
            I => \N__38414\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__38414\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__8051\ : InMux
    port map (
            O => \N__38411\,
            I => \N__38408\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__38408\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__8049\ : CascadeMux
    port map (
            O => \N__38405\,
            I => \N__38402\
        );

    \I__8048\ : InMux
    port map (
            O => \N__38402\,
            I => \N__38399\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__38399\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__8046\ : InMux
    port map (
            O => \N__38396\,
            I => \N__38393\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__38393\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__8044\ : CascadeMux
    port map (
            O => \N__38390\,
            I => \N__38387\
        );

    \I__8043\ : InMux
    port map (
            O => \N__38387\,
            I => \N__38384\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__38384\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__8041\ : InMux
    port map (
            O => \N__38381\,
            I => \N__38378\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__38378\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__8039\ : InMux
    port map (
            O => \N__38375\,
            I => \N__38372\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__38372\,
            I => \N__38368\
        );

    \I__8037\ : InMux
    port map (
            O => \N__38371\,
            I => \N__38365\
        );

    \I__8036\ : Span4Mux_h
    port map (
            O => \N__38368\,
            I => \N__38360\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__38365\,
            I => \N__38360\
        );

    \I__8034\ : Span4Mux_v
    port map (
            O => \N__38360\,
            I => \N__38356\
        );

    \I__8033\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38353\
        );

    \I__8032\ : Odrv4
    port map (
            O => \N__38356\,
            I => measured_delay_tr_10
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__38353\,
            I => measured_delay_tr_10
        );

    \I__8030\ : CascadeMux
    port map (
            O => \N__38348\,
            I => \N__38345\
        );

    \I__8029\ : InMux
    port map (
            O => \N__38345\,
            I => \N__38342\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__38342\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__8027\ : CascadeMux
    port map (
            O => \N__38339\,
            I => \N__38336\
        );

    \I__8026\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38333\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__38333\,
            I => \N__38330\
        );

    \I__8024\ : Odrv4
    port map (
            O => \N__38330\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__8023\ : CascadeMux
    port map (
            O => \N__38327\,
            I => \N__38324\
        );

    \I__8022\ : InMux
    port map (
            O => \N__38324\,
            I => \N__38321\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__38321\,
            I => \N__38318\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__38318\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__38315\,
            I => \N__38308\
        );

    \I__8018\ : InMux
    port map (
            O => \N__38314\,
            I => \N__38298\
        );

    \I__8017\ : InMux
    port map (
            O => \N__38313\,
            I => \N__38298\
        );

    \I__8016\ : InMux
    port map (
            O => \N__38312\,
            I => \N__38298\
        );

    \I__8015\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38298\
        );

    \I__8014\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38292\
        );

    \I__8013\ : InMux
    port map (
            O => \N__38307\,
            I => \N__38292\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__38298\,
            I => \N__38289\
        );

    \I__8011\ : InMux
    port map (
            O => \N__38297\,
            I => \N__38286\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__38292\,
            I => \N__38282\
        );

    \I__8009\ : Span4Mux_h
    port map (
            O => \N__38289\,
            I => \N__38277\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__38286\,
            I => \N__38277\
        );

    \I__8007\ : InMux
    port map (
            O => \N__38285\,
            I => \N__38271\
        );

    \I__8006\ : Span4Mux_v
    port map (
            O => \N__38282\,
            I => \N__38268\
        );

    \I__8005\ : Span4Mux_v
    port map (
            O => \N__38277\,
            I => \N__38265\
        );

    \I__8004\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38258\
        );

    \I__8003\ : InMux
    port map (
            O => \N__38275\,
            I => \N__38258\
        );

    \I__8002\ : InMux
    port map (
            O => \N__38274\,
            I => \N__38258\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__38271\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__8000\ : Odrv4
    port map (
            O => \N__38268\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__7999\ : Odrv4
    port map (
            O => \N__38265\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__38258\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__7997\ : InMux
    port map (
            O => \N__38249\,
            I => \N__38245\
        );

    \I__7996\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38242\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__38245\,
            I => \N__38236\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__38242\,
            I => \N__38236\
        );

    \I__7993\ : InMux
    port map (
            O => \N__38241\,
            I => \N__38233\
        );

    \I__7992\ : Span4Mux_v
    port map (
            O => \N__38236\,
            I => \N__38230\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__38233\,
            I => \N__38227\
        );

    \I__7990\ : Odrv4
    port map (
            O => \N__38230\,
            I => measured_delay_tr_4
        );

    \I__7989\ : Odrv4
    port map (
            O => \N__38227\,
            I => measured_delay_tr_4
        );

    \I__7988\ : CascadeMux
    port map (
            O => \N__38222\,
            I => \N__38219\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38219\,
            I => \N__38216\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__38216\,
            I => \N__38213\
        );

    \I__7985\ : Odrv4
    port map (
            O => \N__38213\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__7984\ : InMux
    port map (
            O => \N__38210\,
            I => \N__38205\
        );

    \I__7983\ : InMux
    port map (
            O => \N__38209\,
            I => \N__38202\
        );

    \I__7982\ : InMux
    port map (
            O => \N__38208\,
            I => \N__38199\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__38205\,
            I => \N__38196\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__38202\,
            I => \N__38193\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__38199\,
            I => \N__38186\
        );

    \I__7978\ : Span4Mux_v
    port map (
            O => \N__38196\,
            I => \N__38186\
        );

    \I__7977\ : Span4Mux_v
    port map (
            O => \N__38193\,
            I => \N__38186\
        );

    \I__7976\ : Odrv4
    port map (
            O => \N__38186\,
            I => \phase_controller_inst2.stoper_tr.time_passed11\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38183\,
            I => \N__38178\
        );

    \I__7974\ : InMux
    port map (
            O => \N__38182\,
            I => \N__38173\
        );

    \I__7973\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38169\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__38178\,
            I => \N__38166\
        );

    \I__7971\ : InMux
    port map (
            O => \N__38177\,
            I => \N__38161\
        );

    \I__7970\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38161\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__38173\,
            I => \N__38158\
        );

    \I__7968\ : InMux
    port map (
            O => \N__38172\,
            I => \N__38155\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__38169\,
            I => \N__38152\
        );

    \I__7966\ : Odrv4
    port map (
            O => \N__38166\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__38161\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7964\ : Odrv4
    port map (
            O => \N__38158\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__38155\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7962\ : Odrv12
    port map (
            O => \N__38152\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7961\ : InMux
    port map (
            O => \N__38141\,
            I => \N__38138\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__38138\,
            I => \N__38135\
        );

    \I__7959\ : Span4Mux_s3_v
    port map (
            O => \N__38135\,
            I => \N__38132\
        );

    \I__7958\ : Odrv4
    port map (
            O => \N__38132\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0\
        );

    \I__7957\ : InMux
    port map (
            O => \N__38129\,
            I => \N__38126\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__38126\,
            I => \N__38123\
        );

    \I__7955\ : Span4Mux_h
    port map (
            O => \N__38123\,
            I => \N__38120\
        );

    \I__7954\ : Odrv4
    port map (
            O => \N__38120\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\
        );

    \I__7953\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38114\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__38114\,
            I => \N__38111\
        );

    \I__7951\ : Span4Mux_v
    port map (
            O => \N__38111\,
            I => \N__38108\
        );

    \I__7950\ : Odrv4
    port map (
            O => \N__38108\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\
        );

    \I__7949\ : CascadeMux
    port map (
            O => \N__38105\,
            I => \N__38102\
        );

    \I__7948\ : InMux
    port map (
            O => \N__38102\,
            I => \N__38088\
        );

    \I__7947\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38081\
        );

    \I__7946\ : InMux
    port map (
            O => \N__38100\,
            I => \N__38081\
        );

    \I__7945\ : InMux
    port map (
            O => \N__38099\,
            I => \N__38081\
        );

    \I__7944\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38078\
        );

    \I__7943\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38069\
        );

    \I__7942\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38069\
        );

    \I__7941\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38069\
        );

    \I__7940\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38069\
        );

    \I__7939\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38060\
        );

    \I__7938\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38060\
        );

    \I__7937\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38060\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__38088\,
            I => \N__38053\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__38081\,
            I => \N__38053\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__38078\,
            I => \N__38053\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__38069\,
            I => \N__38050\
        );

    \I__7932\ : InMux
    port map (
            O => \N__38068\,
            I => \N__38047\
        );

    \I__7931\ : InMux
    port map (
            O => \N__38067\,
            I => \N__38042\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__38060\,
            I => \N__38039\
        );

    \I__7929\ : Sp12to4
    port map (
            O => \N__38053\,
            I => \N__38032\
        );

    \I__7928\ : Sp12to4
    port map (
            O => \N__38050\,
            I => \N__38032\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__38047\,
            I => \N__38032\
        );

    \I__7926\ : InMux
    port map (
            O => \N__38046\,
            I => \N__38027\
        );

    \I__7925\ : InMux
    port map (
            O => \N__38045\,
            I => \N__38027\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__38042\,
            I => \N__38022\
        );

    \I__7923\ : Span4Mux_h
    port map (
            O => \N__38039\,
            I => \N__38022\
        );

    \I__7922\ : Span12Mux_v
    port map (
            O => \N__38032\,
            I => \N__38019\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__38027\,
            I => \N__38014\
        );

    \I__7920\ : Span4Mux_v
    port map (
            O => \N__38022\,
            I => \N__38014\
        );

    \I__7919\ : Odrv12
    port map (
            O => \N__38019\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__7918\ : Odrv4
    port map (
            O => \N__38014\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__7917\ : CascadeMux
    port map (
            O => \N__38009\,
            I => \N__38006\
        );

    \I__7916\ : InMux
    port map (
            O => \N__38006\,
            I => \N__38003\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__38003\,
            I => \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__7914\ : InMux
    port map (
            O => \N__38000\,
            I => \N__37997\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__37997\,
            I => \N__37993\
        );

    \I__7912\ : InMux
    port map (
            O => \N__37996\,
            I => \N__37990\
        );

    \I__7911\ : Sp12to4
    port map (
            O => \N__37993\,
            I => \N__37984\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__37990\,
            I => \N__37984\
        );

    \I__7909\ : InMux
    port map (
            O => \N__37989\,
            I => \N__37981\
        );

    \I__7908\ : Span12Mux_v
    port map (
            O => \N__37984\,
            I => \N__37978\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__37981\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__7906\ : Odrv12
    port map (
            O => \N__37978\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__7905\ : CascadeMux
    port map (
            O => \N__37973\,
            I => \N__37970\
        );

    \I__7904\ : InMux
    port map (
            O => \N__37970\,
            I => \N__37967\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__37967\,
            I => \N__37964\
        );

    \I__7902\ : Odrv12
    port map (
            O => \N__37964\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__7901\ : InMux
    port map (
            O => \N__37961\,
            I => \N__37958\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__37958\,
            I => \N__37954\
        );

    \I__7899\ : InMux
    port map (
            O => \N__37957\,
            I => \N__37951\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__37954\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__37951\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7896\ : InMux
    port map (
            O => \N__37946\,
            I => \N__37943\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__37943\,
            I => \N__37940\
        );

    \I__7894\ : Odrv4
    port map (
            O => \N__37940\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__7893\ : CascadeMux
    port map (
            O => \N__37937\,
            I => \N__37934\
        );

    \I__7892\ : InMux
    port map (
            O => \N__37934\,
            I => \N__37931\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__37931\,
            I => \N__37927\
        );

    \I__7890\ : InMux
    port map (
            O => \N__37930\,
            I => \N__37924\
        );

    \I__7889\ : Odrv4
    port map (
            O => \N__37927\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__37924\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7887\ : InMux
    port map (
            O => \N__37919\,
            I => \N__37916\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__37916\,
            I => \N__37913\
        );

    \I__7885\ : Odrv4
    port map (
            O => \N__37913\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__7884\ : InMux
    port map (
            O => \N__37910\,
            I => \N__37907\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__37907\,
            I => \N__37903\
        );

    \I__7882\ : InMux
    port map (
            O => \N__37906\,
            I => \N__37900\
        );

    \I__7881\ : Odrv12
    port map (
            O => \N__37903\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__37900\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7879\ : CascadeMux
    port map (
            O => \N__37895\,
            I => \N__37892\
        );

    \I__7878\ : InMux
    port map (
            O => \N__37892\,
            I => \N__37889\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__37889\,
            I => \N__37886\
        );

    \I__7876\ : Odrv4
    port map (
            O => \N__37886\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__7875\ : InMux
    port map (
            O => \N__37883\,
            I => \N__37880\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__37880\,
            I => \N__37877\
        );

    \I__7873\ : Span4Mux_s1_v
    port map (
            O => \N__37877\,
            I => \N__37873\
        );

    \I__7872\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37870\
        );

    \I__7871\ : Odrv4
    port map (
            O => \N__37873\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__37870\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7869\ : InMux
    port map (
            O => \N__37865\,
            I => \N__37862\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__37862\,
            I => \N__37859\
        );

    \I__7867\ : Odrv12
    port map (
            O => \N__37859\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__7866\ : InMux
    port map (
            O => \N__37856\,
            I => \N__37853\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__37853\,
            I => \N__37849\
        );

    \I__7864\ : InMux
    port map (
            O => \N__37852\,
            I => \N__37846\
        );

    \I__7863\ : Odrv4
    port map (
            O => \N__37849\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__37846\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7861\ : CascadeMux
    port map (
            O => \N__37841\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__7860\ : CascadeMux
    port map (
            O => \N__37838\,
            I => \N__37835\
        );

    \I__7859\ : InMux
    port map (
            O => \N__37835\,
            I => \N__37831\
        );

    \I__7858\ : InMux
    port map (
            O => \N__37834\,
            I => \N__37827\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__37831\,
            I => \N__37824\
        );

    \I__7856\ : InMux
    port map (
            O => \N__37830\,
            I => \N__37821\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__37827\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7854\ : Odrv12
    port map (
            O => \N__37824\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37821\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7852\ : InMux
    port map (
            O => \N__37814\,
            I => \N__37806\
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__37813\,
            I => \N__37797\
        );

    \I__7850\ : CascadeMux
    port map (
            O => \N__37812\,
            I => \N__37794\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37811\,
            I => \N__37776\
        );

    \I__7848\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37776\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37809\,
            I => \N__37776\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__37806\,
            I => \N__37773\
        );

    \I__7845\ : InMux
    port map (
            O => \N__37805\,
            I => \N__37760\
        );

    \I__7844\ : InMux
    port map (
            O => \N__37804\,
            I => \N__37760\
        );

    \I__7843\ : InMux
    port map (
            O => \N__37803\,
            I => \N__37760\
        );

    \I__7842\ : InMux
    port map (
            O => \N__37802\,
            I => \N__37760\
        );

    \I__7841\ : InMux
    port map (
            O => \N__37801\,
            I => \N__37760\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37800\,
            I => \N__37760\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37797\,
            I => \N__37755\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37755\
        );

    \I__7837\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37746\
        );

    \I__7836\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37746\
        );

    \I__7835\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37746\
        );

    \I__7834\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37746\
        );

    \I__7833\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37739\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37788\,
            I => \N__37739\
        );

    \I__7831\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37739\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37786\,
            I => \N__37734\
        );

    \I__7829\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37734\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__37784\,
            I => \N__37731\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37783\,
            I => \N__37727\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__37776\,
            I => \N__37722\
        );

    \I__7825\ : Span4Mux_v
    port map (
            O => \N__37773\,
            I => \N__37722\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__37760\,
            I => \N__37719\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__37755\,
            I => \N__37710\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__37746\,
            I => \N__37710\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__37739\,
            I => \N__37710\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__37734\,
            I => \N__37710\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37705\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37705\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__37727\,
            I => \N__37702\
        );

    \I__7816\ : Span4Mux_v
    port map (
            O => \N__37722\,
            I => \N__37699\
        );

    \I__7815\ : Span4Mux_h
    port map (
            O => \N__37719\,
            I => \N__37694\
        );

    \I__7814\ : Span4Mux_v
    port map (
            O => \N__37710\,
            I => \N__37694\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__37705\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__7812\ : Odrv4
    port map (
            O => \N__37702\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__37699\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__7810\ : Odrv4
    port map (
            O => \N__37694\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__37685\,
            I => \N__37678\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__37684\,
            I => \N__37668\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37683\,
            I => \N__37656\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37656\
        );

    \I__7805\ : InMux
    port map (
            O => \N__37681\,
            I => \N__37656\
        );

    \I__7804\ : InMux
    port map (
            O => \N__37678\,
            I => \N__37656\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37677\,
            I => \N__37653\
        );

    \I__7802\ : CascadeMux
    port map (
            O => \N__37676\,
            I => \N__37647\
        );

    \I__7801\ : CascadeMux
    port map (
            O => \N__37675\,
            I => \N__37644\
        );

    \I__7800\ : CascadeMux
    port map (
            O => \N__37674\,
            I => \N__37641\
        );

    \I__7799\ : CascadeMux
    port map (
            O => \N__37673\,
            I => \N__37638\
        );

    \I__7798\ : CascadeMux
    port map (
            O => \N__37672\,
            I => \N__37635\
        );

    \I__7797\ : CascadeMux
    port map (
            O => \N__37671\,
            I => \N__37632\
        );

    \I__7796\ : InMux
    port map (
            O => \N__37668\,
            I => \N__37623\
        );

    \I__7795\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37623\
        );

    \I__7794\ : InMux
    port map (
            O => \N__37666\,
            I => \N__37623\
        );

    \I__7793\ : CascadeMux
    port map (
            O => \N__37665\,
            I => \N__37619\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37656\,
            I => \N__37613\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__37653\,
            I => \N__37613\
        );

    \I__7790\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37600\
        );

    \I__7789\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37600\
        );

    \I__7788\ : InMux
    port map (
            O => \N__37650\,
            I => \N__37600\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37647\,
            I => \N__37600\
        );

    \I__7786\ : InMux
    port map (
            O => \N__37644\,
            I => \N__37600\
        );

    \I__7785\ : InMux
    port map (
            O => \N__37641\,
            I => \N__37600\
        );

    \I__7784\ : InMux
    port map (
            O => \N__37638\,
            I => \N__37589\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37635\,
            I => \N__37589\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37632\,
            I => \N__37589\
        );

    \I__7781\ : InMux
    port map (
            O => \N__37631\,
            I => \N__37589\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37630\,
            I => \N__37589\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37623\,
            I => \N__37586\
        );

    \I__7778\ : InMux
    port map (
            O => \N__37622\,
            I => \N__37583\
        );

    \I__7777\ : InMux
    port map (
            O => \N__37619\,
            I => \N__37577\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37618\,
            I => \N__37577\
        );

    \I__7775\ : Span4Mux_s2_v
    port map (
            O => \N__37613\,
            I => \N__37573\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37600\,
            I => \N__37570\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__37589\,
            I => \N__37563\
        );

    \I__7772\ : Span4Mux_v
    port map (
            O => \N__37586\,
            I => \N__37563\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__37583\,
            I => \N__37563\
        );

    \I__7770\ : InMux
    port map (
            O => \N__37582\,
            I => \N__37560\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__37577\,
            I => \N__37557\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37576\,
            I => \N__37554\
        );

    \I__7767\ : Span4Mux_h
    port map (
            O => \N__37573\,
            I => \N__37551\
        );

    \I__7766\ : Span4Mux_h
    port map (
            O => \N__37570\,
            I => \N__37548\
        );

    \I__7765\ : Span4Mux_h
    port map (
            O => \N__37563\,
            I => \N__37545\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__37560\,
            I => \N__37538\
        );

    \I__7763\ : Span4Mux_v
    port map (
            O => \N__37557\,
            I => \N__37538\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__37554\,
            I => \N__37538\
        );

    \I__7761\ : Odrv4
    port map (
            O => \N__37551\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7760\ : Odrv4
    port map (
            O => \N__37548\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7759\ : Odrv4
    port map (
            O => \N__37545\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7758\ : Odrv4
    port map (
            O => \N__37538\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7757\ : CascadeMux
    port map (
            O => \N__37529\,
            I => \N__37519\
        );

    \I__7756\ : InMux
    port map (
            O => \N__37528\,
            I => \N__37500\
        );

    \I__7755\ : InMux
    port map (
            O => \N__37527\,
            I => \N__37500\
        );

    \I__7754\ : InMux
    port map (
            O => \N__37526\,
            I => \N__37500\
        );

    \I__7753\ : InMux
    port map (
            O => \N__37525\,
            I => \N__37500\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37524\,
            I => \N__37500\
        );

    \I__7751\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37497\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__37522\,
            I => \N__37494\
        );

    \I__7749\ : InMux
    port map (
            O => \N__37519\,
            I => \N__37483\
        );

    \I__7748\ : InMux
    port map (
            O => \N__37518\,
            I => \N__37483\
        );

    \I__7747\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37470\
        );

    \I__7746\ : InMux
    port map (
            O => \N__37516\,
            I => \N__37470\
        );

    \I__7745\ : InMux
    port map (
            O => \N__37515\,
            I => \N__37470\
        );

    \I__7744\ : InMux
    port map (
            O => \N__37514\,
            I => \N__37470\
        );

    \I__7743\ : InMux
    port map (
            O => \N__37513\,
            I => \N__37470\
        );

    \I__7742\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37470\
        );

    \I__7741\ : InMux
    port map (
            O => \N__37511\,
            I => \N__37467\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__37500\,
            I => \N__37462\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__37497\,
            I => \N__37462\
        );

    \I__7738\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37457\
        );

    \I__7737\ : InMux
    port map (
            O => \N__37493\,
            I => \N__37457\
        );

    \I__7736\ : InMux
    port map (
            O => \N__37492\,
            I => \N__37454\
        );

    \I__7735\ : InMux
    port map (
            O => \N__37491\,
            I => \N__37445\
        );

    \I__7734\ : InMux
    port map (
            O => \N__37490\,
            I => \N__37445\
        );

    \I__7733\ : InMux
    port map (
            O => \N__37489\,
            I => \N__37445\
        );

    \I__7732\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37445\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__37483\,
            I => \N__37442\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__37470\,
            I => \N__37437\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__37467\,
            I => \N__37432\
        );

    \I__7728\ : Span4Mux_h
    port map (
            O => \N__37462\,
            I => \N__37432\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__37457\,
            I => \N__37427\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__37454\,
            I => \N__37427\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__37445\,
            I => \N__37424\
        );

    \I__7724\ : Span4Mux_s1_v
    port map (
            O => \N__37442\,
            I => \N__37421\
        );

    \I__7723\ : InMux
    port map (
            O => \N__37441\,
            I => \N__37416\
        );

    \I__7722\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37416\
        );

    \I__7721\ : Span4Mux_h
    port map (
            O => \N__37437\,
            I => \N__37413\
        );

    \I__7720\ : Span4Mux_v
    port map (
            O => \N__37432\,
            I => \N__37410\
        );

    \I__7719\ : Span4Mux_h
    port map (
            O => \N__37427\,
            I => \N__37403\
        );

    \I__7718\ : Span4Mux_v
    port map (
            O => \N__37424\,
            I => \N__37403\
        );

    \I__7717\ : Span4Mux_v
    port map (
            O => \N__37421\,
            I => \N__37403\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__37416\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7715\ : Odrv4
    port map (
            O => \N__37413\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7714\ : Odrv4
    port map (
            O => \N__37410\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7713\ : Odrv4
    port map (
            O => \N__37403\,
            I => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7712\ : InMux
    port map (
            O => \N__37394\,
            I => \N__37391\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__37391\,
            I => \N__37388\
        );

    \I__7710\ : Odrv4
    port map (
            O => \N__37388\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__7709\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37382\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__37382\,
            I => \N__37378\
        );

    \I__7707\ : InMux
    port map (
            O => \N__37381\,
            I => \N__37375\
        );

    \I__7706\ : Odrv4
    port map (
            O => \N__37378\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__37375\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7704\ : InMux
    port map (
            O => \N__37370\,
            I => \N__37366\
        );

    \I__7703\ : InMux
    port map (
            O => \N__37369\,
            I => \N__37363\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__37366\,
            I => \N__37360\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__37363\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__7700\ : Odrv12
    port map (
            O => \N__37360\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__7699\ : CascadeMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7698\ : InMux
    port map (
            O => \N__37352\,
            I => \N__37349\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__37349\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__7696\ : InMux
    port map (
            O => \N__37346\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__7695\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37340\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__37340\,
            I => \N__37336\
        );

    \I__7693\ : InMux
    port map (
            O => \N__37339\,
            I => \N__37333\
        );

    \I__7692\ : Span4Mux_v
    port map (
            O => \N__37336\,
            I => \N__37330\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__37333\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__37330\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7689\ : InMux
    port map (
            O => \N__37325\,
            I => \N__37322\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__37322\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__7687\ : InMux
    port map (
            O => \N__37319\,
            I => \bfn_15_4_0_\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37316\,
            I => \N__37312\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37315\,
            I => \N__37309\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__37312\,
            I => \N__37306\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__37309\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7682\ : Odrv12
    port map (
            O => \N__37306\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7681\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37298\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__37298\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__7679\ : InMux
    port map (
            O => \N__37295\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__7678\ : InMux
    port map (
            O => \N__37292\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__7677\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37286\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__37286\,
            I => \N__37283\
        );

    \I__7675\ : Span4Mux_h
    port map (
            O => \N__37283\,
            I => \N__37280\
        );

    \I__7674\ : Odrv4
    port map (
            O => \N__37280\,
            I => \delay_measurement_inst.delay_tr_timer.N_290\
        );

    \I__7673\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37266\
        );

    \I__7672\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37266\
        );

    \I__7671\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37266\
        );

    \I__7670\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37263\
        );

    \I__7669\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37258\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__37266\,
            I => \N__37254\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__37263\,
            I => \N__37251\
        );

    \I__7666\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37246\
        );

    \I__7665\ : InMux
    port map (
            O => \N__37261\,
            I => \N__37246\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__37258\,
            I => \N__37242\
        );

    \I__7663\ : InMux
    port map (
            O => \N__37257\,
            I => \N__37239\
        );

    \I__7662\ : Span4Mux_v
    port map (
            O => \N__37254\,
            I => \N__37232\
        );

    \I__7661\ : Span4Mux_v
    port map (
            O => \N__37251\,
            I => \N__37232\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__37246\,
            I => \N__37232\
        );

    \I__7659\ : InMux
    port map (
            O => \N__37245\,
            I => \N__37229\
        );

    \I__7658\ : Odrv4
    port map (
            O => \N__37242\,
            I => \delay_measurement_inst.N_325\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__37239\,
            I => \delay_measurement_inst.N_325\
        );

    \I__7656\ : Odrv4
    port map (
            O => \N__37232\,
            I => \delay_measurement_inst.N_325\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__37229\,
            I => \delay_measurement_inst.N_325\
        );

    \I__7654\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37217\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__37217\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__7652\ : InMux
    port map (
            O => \N__37214\,
            I => \N__37211\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__37211\,
            I => \N__37207\
        );

    \I__7650\ : InMux
    port map (
            O => \N__37210\,
            I => \N__37204\
        );

    \I__7649\ : Span4Mux_v
    port map (
            O => \N__37207\,
            I => \N__37201\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__37204\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7647\ : Odrv4
    port map (
            O => \N__37201\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7646\ : CascadeMux
    port map (
            O => \N__37196\,
            I => \N__37193\
        );

    \I__7645\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37190\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__37187\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__7642\ : InMux
    port map (
            O => \N__37184\,
            I => \N__37181\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__37181\,
            I => \N__37177\
        );

    \I__7640\ : InMux
    port map (
            O => \N__37180\,
            I => \N__37174\
        );

    \I__7639\ : Odrv4
    port map (
            O => \N__37177\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__37174\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7637\ : InMux
    port map (
            O => \N__37169\,
            I => \N__37166\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__37166\,
            I => \N__37162\
        );

    \I__7635\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37159\
        );

    \I__7634\ : Span4Mux_v
    port map (
            O => \N__37162\,
            I => \N__37156\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__37159\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7632\ : Odrv4
    port map (
            O => \N__37156\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7631\ : InMux
    port map (
            O => \N__37151\,
            I => \N__37148\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__37148\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__7629\ : InMux
    port map (
            O => \N__37145\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__7628\ : InMux
    port map (
            O => \N__37142\,
            I => \N__37138\
        );

    \I__7627\ : InMux
    port map (
            O => \N__37141\,
            I => \N__37135\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__37138\,
            I => \N__37132\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__37135\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7624\ : Odrv4
    port map (
            O => \N__37132\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7623\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__37124\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__7621\ : InMux
    port map (
            O => \N__37121\,
            I => \bfn_15_3_0_\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37118\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__7619\ : InMux
    port map (
            O => \N__37115\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__7618\ : InMux
    port map (
            O => \N__37112\,
            I => \N__37108\
        );

    \I__7617\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37105\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__37108\,
            I => \N__37102\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__37105\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7614\ : Odrv12
    port map (
            O => \N__37102\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__37097\,
            I => \N__37094\
        );

    \I__7612\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37091\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__37091\,
            I => \N__37088\
        );

    \I__7610\ : Odrv12
    port map (
            O => \N__37088\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__7609\ : InMux
    port map (
            O => \N__37085\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__7608\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37078\
        );

    \I__7607\ : InMux
    port map (
            O => \N__37081\,
            I => \N__37075\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__37078\,
            I => \N__37072\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__37075\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7604\ : Odrv12
    port map (
            O => \N__37072\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7603\ : InMux
    port map (
            O => \N__37067\,
            I => \N__37064\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__37064\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__7601\ : InMux
    port map (
            O => \N__37061\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__7600\ : InMux
    port map (
            O => \N__37058\,
            I => \N__37054\
        );

    \I__7599\ : InMux
    port map (
            O => \N__37057\,
            I => \N__37051\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__37054\,
            I => \N__37048\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__37051\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7596\ : Odrv4
    port map (
            O => \N__37048\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7595\ : InMux
    port map (
            O => \N__37043\,
            I => \N__37040\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__37040\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__7593\ : InMux
    port map (
            O => \N__37037\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__7592\ : InMux
    port map (
            O => \N__37034\,
            I => \N__37031\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__37031\,
            I => \N__37027\
        );

    \I__7590\ : InMux
    port map (
            O => \N__37030\,
            I => \N__37024\
        );

    \I__7589\ : Span4Mux_v
    port map (
            O => \N__37027\,
            I => \N__37021\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__37024\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7587\ : Odrv4
    port map (
            O => \N__37021\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7586\ : CascadeMux
    port map (
            O => \N__37016\,
            I => \N__37013\
        );

    \I__7585\ : InMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__37010\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__7583\ : InMux
    port map (
            O => \N__37007\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__7582\ : InMux
    port map (
            O => \N__37004\,
            I => \N__36998\
        );

    \I__7581\ : InMux
    port map (
            O => \N__37003\,
            I => \N__36993\
        );

    \I__7580\ : InMux
    port map (
            O => \N__37002\,
            I => \N__36993\
        );

    \I__7579\ : InMux
    port map (
            O => \N__37001\,
            I => \N__36990\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__36998\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__36993\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__36990\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7575\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36975\
        );

    \I__7574\ : InMux
    port map (
            O => \N__36982\,
            I => \N__36975\
        );

    \I__7573\ : InMux
    port map (
            O => \N__36981\,
            I => \N__36972\
        );

    \I__7572\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36969\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__36975\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__36972\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__36969\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7568\ : InMux
    port map (
            O => \N__36962\,
            I => \N__36959\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__36959\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__7566\ : InMux
    port map (
            O => \N__36956\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__7565\ : InMux
    port map (
            O => \N__36953\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__7564\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36946\
        );

    \I__7563\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36943\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__36946\,
            I => \N__36940\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__36943\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__36940\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7559\ : InMux
    port map (
            O => \N__36935\,
            I => \N__36932\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__36932\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__7557\ : InMux
    port map (
            O => \N__36929\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__7556\ : InMux
    port map (
            O => \N__36926\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__7555\ : InMux
    port map (
            O => \N__36923\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__7554\ : InMux
    port map (
            O => \N__36920\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__7553\ : InMux
    port map (
            O => \N__36917\,
            I => \N__36913\
        );

    \I__7552\ : InMux
    port map (
            O => \N__36916\,
            I => \N__36910\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__36913\,
            I => \N__36907\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__36910\,
            I => \N__36904\
        );

    \I__7549\ : Span4Mux_v
    port map (
            O => \N__36907\,
            I => \N__36900\
        );

    \I__7548\ : Span4Mux_h
    port map (
            O => \N__36904\,
            I => \N__36897\
        );

    \I__7547\ : InMux
    port map (
            O => \N__36903\,
            I => \N__36894\
        );

    \I__7546\ : Odrv4
    port map (
            O => \N__36900\,
            I => \phase_controller_inst2.stoper_hc.time_passed11\
        );

    \I__7545\ : Odrv4
    port map (
            O => \N__36897\,
            I => \phase_controller_inst2.stoper_hc.time_passed11\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__36894\,
            I => \phase_controller_inst2.stoper_hc.time_passed11\
        );

    \I__7543\ : CascadeMux
    port map (
            O => \N__36887\,
            I => \N__36884\
        );

    \I__7542\ : InMux
    port map (
            O => \N__36884\,
            I => \N__36881\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__36881\,
            I => \N__36878\
        );

    \I__7540\ : Span4Mux_v
    port map (
            O => \N__36878\,
            I => \N__36875\
        );

    \I__7539\ : Odrv4
    port map (
            O => \N__36875\,
            I => \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__7538\ : CascadeMux
    port map (
            O => \N__36872\,
            I => \N__36869\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36865\
        );

    \I__7536\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36862\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__36865\,
            I => \N__36857\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36854\
        );

    \I__7533\ : InMux
    port map (
            O => \N__36861\,
            I => \N__36851\
        );

    \I__7532\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36846\
        );

    \I__7531\ : Span4Mux_v
    port map (
            O => \N__36857\,
            I => \N__36843\
        );

    \I__7530\ : Span4Mux_v
    port map (
            O => \N__36854\,
            I => \N__36840\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__36851\,
            I => \N__36837\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36850\,
            I => \N__36834\
        );

    \I__7527\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36831\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__36846\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7525\ : Odrv4
    port map (
            O => \N__36843\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7524\ : Odrv4
    port map (
            O => \N__36840\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7523\ : Odrv4
    port map (
            O => \N__36837\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__36834\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__36831\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7520\ : InMux
    port map (
            O => \N__36818\,
            I => \N__36815\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__36815\,
            I => \N__36812\
        );

    \I__7518\ : Span4Mux_h
    port map (
            O => \N__36812\,
            I => \N__36809\
        );

    \I__7517\ : Span4Mux_h
    port map (
            O => \N__36809\,
            I => \N__36803\
        );

    \I__7516\ : InMux
    port map (
            O => \N__36808\,
            I => \N__36798\
        );

    \I__7515\ : InMux
    port map (
            O => \N__36807\,
            I => \N__36798\
        );

    \I__7514\ : InMux
    port map (
            O => \N__36806\,
            I => \N__36795\
        );

    \I__7513\ : Sp12to4
    port map (
            O => \N__36803\,
            I => \N__36790\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__36798\,
            I => \N__36790\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__36795\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__7510\ : Odrv12
    port map (
            O => \N__36790\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__7509\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36782\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__36782\,
            I => \N__36779\
        );

    \I__7507\ : Odrv12
    port map (
            O => \N__36779\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__7506\ : InMux
    port map (
            O => \N__36776\,
            I => \N__36773\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__36773\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__7504\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36767\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__7502\ : Span12Mux_v
    port map (
            O => \N__36764\,
            I => \N__36761\
        );

    \I__7501\ : Odrv12
    port map (
            O => \N__36761\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36758\,
            I => \N__36755\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__36755\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__7498\ : InMux
    port map (
            O => \N__36752\,
            I => \N__36749\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__36749\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__7496\ : CascadeMux
    port map (
            O => \N__36746\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__7495\ : InMux
    port map (
            O => \N__36743\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__7494\ : InMux
    port map (
            O => \N__36740\,
            I => \N__36737\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__36737\,
            I => \N__36734\
        );

    \I__7492\ : Span12Mux_h
    port map (
            O => \N__36734\,
            I => \N__36731\
        );

    \I__7491\ : Odrv12
    port map (
            O => \N__36731\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__7490\ : InMux
    port map (
            O => \N__36728\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36722\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__36722\,
            I => \N__36719\
        );

    \I__7487\ : Span4Mux_h
    port map (
            O => \N__36719\,
            I => \N__36716\
        );

    \I__7486\ : Span4Mux_v
    port map (
            O => \N__36716\,
            I => \N__36713\
        );

    \I__7485\ : Span4Mux_h
    port map (
            O => \N__36713\,
            I => \N__36710\
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__36710\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__7483\ : InMux
    port map (
            O => \N__36707\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__7482\ : InMux
    port map (
            O => \N__36704\,
            I => \N__36701\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__36701\,
            I => \N__36698\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__36698\,
            I => \N__36695\
        );

    \I__7479\ : Odrv4
    port map (
            O => \N__36695\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36692\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36689\,
            I => \N__36686\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__36686\,
            I => \N__36683\
        );

    \I__7475\ : Span4Mux_h
    port map (
            O => \N__36683\,
            I => \N__36680\
        );

    \I__7474\ : Span4Mux_v
    port map (
            O => \N__36680\,
            I => \N__36677\
        );

    \I__7473\ : Span4Mux_h
    port map (
            O => \N__36677\,
            I => \N__36674\
        );

    \I__7472\ : Odrv4
    port map (
            O => \N__36674\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__7471\ : InMux
    port map (
            O => \N__36671\,
            I => \bfn_14_17_0_\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36668\,
            I => \N__36665\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__36665\,
            I => \N__36662\
        );

    \I__7468\ : Odrv4
    port map (
            O => \N__36662\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__7467\ : InMux
    port map (
            O => \N__36659\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__7466\ : InMux
    port map (
            O => \N__36656\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__7465\ : InMux
    port map (
            O => \N__36653\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__7464\ : InMux
    port map (
            O => \N__36650\,
            I => \N__36647\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__36647\,
            I => \N__36643\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36640\
        );

    \I__7461\ : Span4Mux_v
    port map (
            O => \N__36643\,
            I => \N__36635\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__36640\,
            I => \N__36635\
        );

    \I__7459\ : Span4Mux_v
    port map (
            O => \N__36635\,
            I => \N__36632\
        );

    \I__7458\ : Odrv4
    port map (
            O => \N__36632\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__7457\ : CascadeMux
    port map (
            O => \N__36629\,
            I => \N__36623\
        );

    \I__7456\ : CascadeMux
    port map (
            O => \N__36628\,
            I => \N__36616\
        );

    \I__7455\ : CascadeMux
    port map (
            O => \N__36627\,
            I => \N__36613\
        );

    \I__7454\ : CascadeMux
    port map (
            O => \N__36626\,
            I => \N__36610\
        );

    \I__7453\ : InMux
    port map (
            O => \N__36623\,
            I => \N__36598\
        );

    \I__7452\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36583\
        );

    \I__7451\ : InMux
    port map (
            O => \N__36621\,
            I => \N__36583\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36620\,
            I => \N__36583\
        );

    \I__7449\ : InMux
    port map (
            O => \N__36619\,
            I => \N__36583\
        );

    \I__7448\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36583\
        );

    \I__7447\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36583\
        );

    \I__7446\ : InMux
    port map (
            O => \N__36610\,
            I => \N__36583\
        );

    \I__7445\ : CascadeMux
    port map (
            O => \N__36609\,
            I => \N__36580\
        );

    \I__7444\ : InMux
    port map (
            O => \N__36608\,
            I => \N__36576\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36607\,
            I => \N__36573\
        );

    \I__7442\ : InMux
    port map (
            O => \N__36606\,
            I => \N__36570\
        );

    \I__7441\ : CascadeMux
    port map (
            O => \N__36605\,
            I => \N__36567\
        );

    \I__7440\ : CascadeMux
    port map (
            O => \N__36604\,
            I => \N__36563\
        );

    \I__7439\ : CascadeMux
    port map (
            O => \N__36603\,
            I => \N__36560\
        );

    \I__7438\ : CascadeMux
    port map (
            O => \N__36602\,
            I => \N__36557\
        );

    \I__7437\ : CascadeMux
    port map (
            O => \N__36601\,
            I => \N__36554\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36598\,
            I => \N__36544\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__36583\,
            I => \N__36544\
        );

    \I__7434\ : InMux
    port map (
            O => \N__36580\,
            I => \N__36539\
        );

    \I__7433\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36539\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__36576\,
            I => \N__36536\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__36573\,
            I => \N__36533\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36570\,
            I => \N__36530\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36567\,
            I => \N__36527\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36566\,
            I => \N__36510\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36510\
        );

    \I__7426\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36510\
        );

    \I__7425\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36510\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36510\
        );

    \I__7423\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36510\
        );

    \I__7422\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36510\
        );

    \I__7421\ : InMux
    port map (
            O => \N__36551\,
            I => \N__36510\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36550\,
            I => \N__36505\
        );

    \I__7419\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36505\
        );

    \I__7418\ : Span4Mux_v
    port map (
            O => \N__36544\,
            I => \N__36502\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__36539\,
            I => \N__36493\
        );

    \I__7416\ : Span4Mux_v
    port map (
            O => \N__36536\,
            I => \N__36493\
        );

    \I__7415\ : Span4Mux_v
    port map (
            O => \N__36533\,
            I => \N__36493\
        );

    \I__7414\ : Span4Mux_h
    port map (
            O => \N__36530\,
            I => \N__36493\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__36527\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__36510\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__36505\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__7410\ : Odrv4
    port map (
            O => \N__36502\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__36493\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__7408\ : CascadeMux
    port map (
            O => \N__36482\,
            I => \N__36460\
        );

    \I__7407\ : CascadeMux
    port map (
            O => \N__36481\,
            I => \N__36456\
        );

    \I__7406\ : CascadeMux
    port map (
            O => \N__36480\,
            I => \N__36453\
        );

    \I__7405\ : CascadeMux
    port map (
            O => \N__36479\,
            I => \N__36450\
        );

    \I__7404\ : CascadeMux
    port map (
            O => \N__36478\,
            I => \N__36447\
        );

    \I__7403\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36443\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36476\,
            I => \N__36440\
        );

    \I__7401\ : InMux
    port map (
            O => \N__36475\,
            I => \N__36431\
        );

    \I__7400\ : InMux
    port map (
            O => \N__36474\,
            I => \N__36431\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36473\,
            I => \N__36431\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36472\,
            I => \N__36431\
        );

    \I__7397\ : InMux
    port map (
            O => \N__36471\,
            I => \N__36428\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36470\,
            I => \N__36412\
        );

    \I__7395\ : InMux
    port map (
            O => \N__36469\,
            I => \N__36412\
        );

    \I__7394\ : InMux
    port map (
            O => \N__36468\,
            I => \N__36412\
        );

    \I__7393\ : InMux
    port map (
            O => \N__36467\,
            I => \N__36412\
        );

    \I__7392\ : InMux
    port map (
            O => \N__36466\,
            I => \N__36412\
        );

    \I__7391\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36412\
        );

    \I__7390\ : InMux
    port map (
            O => \N__36464\,
            I => \N__36412\
        );

    \I__7389\ : InMux
    port map (
            O => \N__36463\,
            I => \N__36409\
        );

    \I__7388\ : InMux
    port map (
            O => \N__36460\,
            I => \N__36406\
        );

    \I__7387\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36403\
        );

    \I__7386\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36394\
        );

    \I__7385\ : InMux
    port map (
            O => \N__36453\,
            I => \N__36394\
        );

    \I__7384\ : InMux
    port map (
            O => \N__36450\,
            I => \N__36394\
        );

    \I__7383\ : InMux
    port map (
            O => \N__36447\,
            I => \N__36394\
        );

    \I__7382\ : InMux
    port map (
            O => \N__36446\,
            I => \N__36391\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__36443\,
            I => \N__36388\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__36440\,
            I => \N__36385\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__36431\,
            I => \N__36380\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__36428\,
            I => \N__36380\
        );

    \I__7377\ : InMux
    port map (
            O => \N__36427\,
            I => \N__36377\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__36412\,
            I => \N__36373\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__36409\,
            I => \N__36366\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__36406\,
            I => \N__36366\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__36403\,
            I => \N__36366\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__36394\,
            I => \N__36353\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__36391\,
            I => \N__36353\
        );

    \I__7370\ : Span4Mux_h
    port map (
            O => \N__36388\,
            I => \N__36353\
        );

    \I__7369\ : Span4Mux_v
    port map (
            O => \N__36385\,
            I => \N__36353\
        );

    \I__7368\ : Span4Mux_h
    port map (
            O => \N__36380\,
            I => \N__36353\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__36377\,
            I => \N__36353\
        );

    \I__7366\ : InMux
    port map (
            O => \N__36376\,
            I => \N__36350\
        );

    \I__7365\ : Span4Mux_v
    port map (
            O => \N__36373\,
            I => \N__36347\
        );

    \I__7364\ : Span4Mux_v
    port map (
            O => \N__36366\,
            I => \N__36344\
        );

    \I__7363\ : Span4Mux_v
    port map (
            O => \N__36353\,
            I => \N__36341\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__36350\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__7361\ : Odrv4
    port map (
            O => \N__36347\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__7360\ : Odrv4
    port map (
            O => \N__36344\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__36341\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__7358\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36312\
        );

    \I__7357\ : InMux
    port map (
            O => \N__36331\,
            I => \N__36297\
        );

    \I__7356\ : InMux
    port map (
            O => \N__36330\,
            I => \N__36297\
        );

    \I__7355\ : InMux
    port map (
            O => \N__36329\,
            I => \N__36297\
        );

    \I__7354\ : InMux
    port map (
            O => \N__36328\,
            I => \N__36297\
        );

    \I__7353\ : InMux
    port map (
            O => \N__36327\,
            I => \N__36297\
        );

    \I__7352\ : InMux
    port map (
            O => \N__36326\,
            I => \N__36297\
        );

    \I__7351\ : InMux
    port map (
            O => \N__36325\,
            I => \N__36297\
        );

    \I__7350\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36293\
        );

    \I__7349\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36290\
        );

    \I__7348\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36270\
        );

    \I__7347\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36270\
        );

    \I__7346\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36270\
        );

    \I__7345\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36270\
        );

    \I__7344\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36270\
        );

    \I__7343\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36270\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36270\
        );

    \I__7341\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36270\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__36312\,
            I => \N__36267\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__36297\,
            I => \N__36264\
        );

    \I__7338\ : InMux
    port map (
            O => \N__36296\,
            I => \N__36261\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__36293\,
            I => \N__36258\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__36290\,
            I => \N__36255\
        );

    \I__7335\ : InMux
    port map (
            O => \N__36289\,
            I => \N__36250\
        );

    \I__7334\ : InMux
    port map (
            O => \N__36288\,
            I => \N__36245\
        );

    \I__7333\ : InMux
    port map (
            O => \N__36287\,
            I => \N__36245\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__36270\,
            I => \N__36238\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__36267\,
            I => \N__36238\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__36264\,
            I => \N__36238\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__36261\,
            I => \N__36235\
        );

    \I__7328\ : Span4Mux_h
    port map (
            O => \N__36258\,
            I => \N__36230\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__36255\,
            I => \N__36230\
        );

    \I__7326\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36225\
        );

    \I__7325\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36225\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__36250\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__36245\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__7322\ : Odrv4
    port map (
            O => \N__36238\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__7321\ : Odrv12
    port map (
            O => \N__36235\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__36230\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__36225\,
            I => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__7318\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36209\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__36209\,
            I => \N__36202\
        );

    \I__7316\ : InMux
    port map (
            O => \N__36208\,
            I => \N__36199\
        );

    \I__7315\ : CascadeMux
    port map (
            O => \N__36207\,
            I => \N__36196\
        );

    \I__7314\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36193\
        );

    \I__7313\ : CascadeMux
    port map (
            O => \N__36205\,
            I => \N__36190\
        );

    \I__7312\ : Span4Mux_v
    port map (
            O => \N__36202\,
            I => \N__36187\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__36199\,
            I => \N__36184\
        );

    \I__7310\ : InMux
    port map (
            O => \N__36196\,
            I => \N__36181\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__36193\,
            I => \N__36178\
        );

    \I__7308\ : InMux
    port map (
            O => \N__36190\,
            I => \N__36175\
        );

    \I__7307\ : Span4Mux_v
    port map (
            O => \N__36187\,
            I => \N__36172\
        );

    \I__7306\ : Span4Mux_h
    port map (
            O => \N__36184\,
            I => \N__36169\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__36181\,
            I => \N__36164\
        );

    \I__7304\ : Span4Mux_h
    port map (
            O => \N__36178\,
            I => \N__36164\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__36175\,
            I => measured_delay_hc_31
        );

    \I__7302\ : Odrv4
    port map (
            O => \N__36172\,
            I => measured_delay_hc_31
        );

    \I__7301\ : Odrv4
    port map (
            O => \N__36169\,
            I => measured_delay_hc_31
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__36164\,
            I => measured_delay_hc_31
        );

    \I__7299\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36152\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__36152\,
            I => \N__36149\
        );

    \I__7297\ : Span4Mux_h
    port map (
            O => \N__36149\,
            I => \N__36144\
        );

    \I__7296\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36141\
        );

    \I__7295\ : InMux
    port map (
            O => \N__36147\,
            I => \N__36138\
        );

    \I__7294\ : Odrv4
    port map (
            O => \N__36144\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__36141\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__36138\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__7291\ : InMux
    port map (
            O => \N__36131\,
            I => \N__36127\
        );

    \I__7290\ : InMux
    port map (
            O => \N__36130\,
            I => \N__36124\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__36127\,
            I => \N__36117\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__36124\,
            I => \N__36117\
        );

    \I__7287\ : InMux
    port map (
            O => \N__36123\,
            I => \N__36114\
        );

    \I__7286\ : InMux
    port map (
            O => \N__36122\,
            I => \N__36111\
        );

    \I__7285\ : Span4Mux_v
    port map (
            O => \N__36117\,
            I => \N__36108\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__36114\,
            I => \N__36105\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__36111\,
            I => \N__36102\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__36108\,
            I => \N__36099\
        );

    \I__7281\ : Span4Mux_h
    port map (
            O => \N__36105\,
            I => \N__36096\
        );

    \I__7280\ : Odrv12
    port map (
            O => \N__36102\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1\
        );

    \I__7279\ : Odrv4
    port map (
            O => \N__36099\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1\
        );

    \I__7278\ : Odrv4
    port map (
            O => \N__36096\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1\
        );

    \I__7277\ : CascadeMux
    port map (
            O => \N__36089\,
            I => \N__36086\
        );

    \I__7276\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36083\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__36083\,
            I => \N__36080\
        );

    \I__7274\ : Odrv4
    port map (
            O => \N__36080\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__7273\ : CEMux
    port map (
            O => \N__36077\,
            I => \N__36072\
        );

    \I__7272\ : CEMux
    port map (
            O => \N__36076\,
            I => \N__36069\
        );

    \I__7271\ : CEMux
    port map (
            O => \N__36075\,
            I => \N__36066\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__36072\,
            I => \N__36063\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__36069\,
            I => \N__36059\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__36066\,
            I => \N__36056\
        );

    \I__7267\ : Span4Mux_v
    port map (
            O => \N__36063\,
            I => \N__36053\
        );

    \I__7266\ : CEMux
    port map (
            O => \N__36062\,
            I => \N__36050\
        );

    \I__7265\ : Span4Mux_v
    port map (
            O => \N__36059\,
            I => \N__36047\
        );

    \I__7264\ : Span4Mux_h
    port map (
            O => \N__36056\,
            I => \N__36044\
        );

    \I__7263\ : Sp12to4
    port map (
            O => \N__36053\,
            I => \N__36039\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__36050\,
            I => \N__36039\
        );

    \I__7261\ : Span4Mux_h
    port map (
            O => \N__36047\,
            I => \N__36036\
        );

    \I__7260\ : Odrv4
    port map (
            O => \N__36044\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__7259\ : Odrv12
    port map (
            O => \N__36039\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__36036\,
            I => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__7257\ : CascadeMux
    port map (
            O => \N__36029\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__7256\ : InMux
    port map (
            O => \N__36026\,
            I => \N__36023\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__36023\,
            I => \N__36020\
        );

    \I__7254\ : Span4Mux_h
    port map (
            O => \N__36020\,
            I => \N__36017\
        );

    \I__7253\ : Odrv4
    port map (
            O => \N__36017\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0\
        );

    \I__7252\ : InMux
    port map (
            O => \N__36014\,
            I => \N__36010\
        );

    \I__7251\ : InMux
    port map (
            O => \N__36013\,
            I => \N__36007\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__36010\,
            I => \N__36004\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__36007\,
            I => \N__36001\
        );

    \I__7248\ : Span4Mux_v
    port map (
            O => \N__36004\,
            I => \N__35998\
        );

    \I__7247\ : Span12Mux_v
    port map (
            O => \N__36001\,
            I => \N__35995\
        );

    \I__7246\ : Span4Mux_v
    port map (
            O => \N__35998\,
            I => \N__35992\
        );

    \I__7245\ : Odrv12
    port map (
            O => \N__35995\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__7244\ : Odrv4
    port map (
            O => \N__35992\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__7243\ : InMux
    port map (
            O => \N__35987\,
            I => \N__35984\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__35984\,
            I => \N__35981\
        );

    \I__7241\ : Span4Mux_v
    port map (
            O => \N__35981\,
            I => \N__35978\
        );

    \I__7240\ : Odrv4
    port map (
            O => \N__35978\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__7239\ : InMux
    port map (
            O => \N__35975\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__7238\ : InMux
    port map (
            O => \N__35972\,
            I => \N__35969\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__35969\,
            I => \N__35966\
        );

    \I__7236\ : Span4Mux_h
    port map (
            O => \N__35966\,
            I => \N__35963\
        );

    \I__7235\ : Span4Mux_v
    port map (
            O => \N__35963\,
            I => \N__35960\
        );

    \I__7234\ : Span4Mux_h
    port map (
            O => \N__35960\,
            I => \N__35957\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__35957\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35954\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__7231\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35948\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__35948\,
            I => \N__35945\
        );

    \I__7229\ : Span4Mux_v
    port map (
            O => \N__35945\,
            I => \N__35942\
        );

    \I__7228\ : Odrv4
    port map (
            O => \N__35942\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__7227\ : InMux
    port map (
            O => \N__35939\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__7226\ : InMux
    port map (
            O => \N__35936\,
            I => \N__35933\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__35933\,
            I => \N__35930\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__35930\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__7223\ : CEMux
    port map (
            O => \N__35927\,
            I => \N__35924\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__35924\,
            I => \N__35921\
        );

    \I__7221\ : Span4Mux_v
    port map (
            O => \N__35921\,
            I => \N__35917\
        );

    \I__7220\ : CEMux
    port map (
            O => \N__35920\,
            I => \N__35914\
        );

    \I__7219\ : Span4Mux_v
    port map (
            O => \N__35917\,
            I => \N__35908\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__35914\,
            I => \N__35908\
        );

    \I__7217\ : IoInMux
    port map (
            O => \N__35913\,
            I => \N__35905\
        );

    \I__7216\ : Span4Mux_h
    port map (
            O => \N__35908\,
            I => \N__35901\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__35905\,
            I => \N__35897\
        );

    \I__7214\ : CEMux
    port map (
            O => \N__35904\,
            I => \N__35894\
        );

    \I__7213\ : Span4Mux_v
    port map (
            O => \N__35901\,
            I => \N__35891\
        );

    \I__7212\ : CEMux
    port map (
            O => \N__35900\,
            I => \N__35888\
        );

    \I__7211\ : Span4Mux_s1_v
    port map (
            O => \N__35897\,
            I => \N__35885\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__35894\,
            I => \N__35882\
        );

    \I__7209\ : Span4Mux_v
    port map (
            O => \N__35891\,
            I => \N__35877\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__35888\,
            I => \N__35877\
        );

    \I__7207\ : Sp12to4
    port map (
            O => \N__35885\,
            I => \N__35874\
        );

    \I__7206\ : Span4Mux_v
    port map (
            O => \N__35882\,
            I => \N__35871\
        );

    \I__7205\ : Span4Mux_h
    port map (
            O => \N__35877\,
            I => \N__35868\
        );

    \I__7204\ : Span12Mux_h
    port map (
            O => \N__35874\,
            I => \N__35865\
        );

    \I__7203\ : Span4Mux_v
    port map (
            O => \N__35871\,
            I => \N__35862\
        );

    \I__7202\ : Span4Mux_v
    port map (
            O => \N__35868\,
            I => \N__35859\
        );

    \I__7201\ : Span12Mux_v
    port map (
            O => \N__35865\,
            I => \N__35856\
        );

    \I__7200\ : Span4Mux_v
    port map (
            O => \N__35862\,
            I => \N__35853\
        );

    \I__7199\ : Span4Mux_v
    port map (
            O => \N__35859\,
            I => \N__35850\
        );

    \I__7198\ : Odrv12
    port map (
            O => \N__35856\,
            I => red_c_i
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__35853\,
            I => red_c_i
        );

    \I__7196\ : Odrv4
    port map (
            O => \N__35850\,
            I => red_c_i
        );

    \I__7195\ : InMux
    port map (
            O => \N__35843\,
            I => \N__35840\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__35840\,
            I => \N__35837\
        );

    \I__7193\ : Odrv4
    port map (
            O => \N__35837\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__7192\ : CascadeMux
    port map (
            O => \N__35834\,
            I => \phase_controller_inst2.start_timer_hc_RNO_0_0_cascade_\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35831\,
            I => \N__35828\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__35828\,
            I => \N__35823\
        );

    \I__7189\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35819\
        );

    \I__7188\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35816\
        );

    \I__7187\ : Span4Mux_v
    port map (
            O => \N__35823\,
            I => \N__35813\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__35822\,
            I => \N__35810\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__35819\,
            I => \N__35805\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__35816\,
            I => \N__35805\
        );

    \I__7183\ : Span4Mux_v
    port map (
            O => \N__35813\,
            I => \N__35802\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35799\
        );

    \I__7181\ : Span4Mux_h
    port map (
            O => \N__35805\,
            I => \N__35796\
        );

    \I__7180\ : Odrv4
    port map (
            O => \N__35802\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__35799\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__35796\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35789\,
            I => \N__35786\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__35786\,
            I => \N__35782\
        );

    \I__7175\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35778\
        );

    \I__7174\ : Span4Mux_v
    port map (
            O => \N__35782\,
            I => \N__35775\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35772\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__35778\,
            I => \N__35765\
        );

    \I__7171\ : Sp12to4
    port map (
            O => \N__35775\,
            I => \N__35765\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__35772\,
            I => \N__35765\
        );

    \I__7169\ : Odrv12
    port map (
            O => \N__35765\,
            I => \il_max_comp2_D2\
        );

    \I__7168\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35759\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__35759\,
            I => \N__35756\
        );

    \I__7166\ : Span4Mux_h
    port map (
            O => \N__35756\,
            I => \N__35753\
        );

    \I__7165\ : Span4Mux_h
    port map (
            O => \N__35753\,
            I => \N__35749\
        );

    \I__7164\ : CascadeMux
    port map (
            O => \N__35752\,
            I => \N__35746\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__35749\,
            I => \N__35742\
        );

    \I__7162\ : InMux
    port map (
            O => \N__35746\,
            I => \N__35737\
        );

    \I__7161\ : InMux
    port map (
            O => \N__35745\,
            I => \N__35737\
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__35742\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__35737\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__7158\ : InMux
    port map (
            O => \N__35732\,
            I => \N__35729\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35729\,
            I => \N__35726\
        );

    \I__7156\ : Odrv4
    port map (
            O => \N__35726\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35720\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__35720\,
            I => \N__35716\
        );

    \I__7153\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35713\
        );

    \I__7152\ : Odrv4
    port map (
            O => \N__35716\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__35713\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7150\ : CascadeMux
    port map (
            O => \N__35708\,
            I => \phase_controller_inst2.stoper_hc.time_passed11_cascade_\
        );

    \I__7149\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35702\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__35702\,
            I => \N__35699\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__35699\,
            I => \N__35696\
        );

    \I__7146\ : Odrv4
    port map (
            O => \N__35696\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__7145\ : CascadeMux
    port map (
            O => \N__35693\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__7144\ : CascadeMux
    port map (
            O => \N__35690\,
            I => \N__35687\
        );

    \I__7143\ : InMux
    port map (
            O => \N__35687\,
            I => \N__35684\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__35684\,
            I => \N__35680\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35676\
        );

    \I__7140\ : Span4Mux_v
    port map (
            O => \N__35680\,
            I => \N__35673\
        );

    \I__7139\ : InMux
    port map (
            O => \N__35679\,
            I => \N__35670\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__35676\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__35673\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__35670\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7135\ : InMux
    port map (
            O => \N__35663\,
            I => \N__35660\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__35660\,
            I => \N__35657\
        );

    \I__7133\ : Span4Mux_h
    port map (
            O => \N__35657\,
            I => \N__35654\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__35654\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__7131\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35648\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35648\,
            I => \N__35645\
        );

    \I__7129\ : Span4Mux_h
    port map (
            O => \N__35645\,
            I => \N__35641\
        );

    \I__7128\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35638\
        );

    \I__7127\ : Odrv4
    port map (
            O => \N__35641\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__35638\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35626\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35626\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35623\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__35626\,
            I => \N__35620\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__35623\,
            I => \N__35616\
        );

    \I__7120\ : Span4Mux_v
    port map (
            O => \N__35620\,
            I => \N__35613\
        );

    \I__7119\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35610\
        );

    \I__7118\ : Span4Mux_v
    port map (
            O => \N__35616\,
            I => \N__35602\
        );

    \I__7117\ : Span4Mux_h
    port map (
            O => \N__35613\,
            I => \N__35602\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__35610\,
            I => \N__35602\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35598\
        );

    \I__7114\ : Span4Mux_h
    port map (
            O => \N__35602\,
            I => \N__35595\
        );

    \I__7113\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35592\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__35598\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7111\ : Odrv4
    port map (
            O => \N__35595\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35592\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__7109\ : CascadeMux
    port map (
            O => \N__35585\,
            I => \N__35575\
        );

    \I__7108\ : CascadeMux
    port map (
            O => \N__35584\,
            I => \N__35568\
        );

    \I__7107\ : CascadeMux
    port map (
            O => \N__35583\,
            I => \N__35565\
        );

    \I__7106\ : CascadeMux
    port map (
            O => \N__35582\,
            I => \N__35562\
        );

    \I__7105\ : CascadeMux
    port map (
            O => \N__35581\,
            I => \N__35559\
        );

    \I__7104\ : CascadeMux
    port map (
            O => \N__35580\,
            I => \N__35556\
        );

    \I__7103\ : CascadeMux
    port map (
            O => \N__35579\,
            I => \N__35553\
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__35578\,
            I => \N__35550\
        );

    \I__7101\ : InMux
    port map (
            O => \N__35575\,
            I => \N__35537\
        );

    \I__7100\ : InMux
    port map (
            O => \N__35574\,
            I => \N__35537\
        );

    \I__7099\ : CascadeMux
    port map (
            O => \N__35573\,
            I => \N__35534\
        );

    \I__7098\ : CascadeMux
    port map (
            O => \N__35572\,
            I => \N__35531\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__35571\,
            I => \N__35528\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35520\
        );

    \I__7095\ : InMux
    port map (
            O => \N__35565\,
            I => \N__35520\
        );

    \I__7094\ : InMux
    port map (
            O => \N__35562\,
            I => \N__35520\
        );

    \I__7093\ : InMux
    port map (
            O => \N__35559\,
            I => \N__35503\
        );

    \I__7092\ : InMux
    port map (
            O => \N__35556\,
            I => \N__35503\
        );

    \I__7091\ : InMux
    port map (
            O => \N__35553\,
            I => \N__35503\
        );

    \I__7090\ : InMux
    port map (
            O => \N__35550\,
            I => \N__35503\
        );

    \I__7089\ : InMux
    port map (
            O => \N__35549\,
            I => \N__35503\
        );

    \I__7088\ : InMux
    port map (
            O => \N__35548\,
            I => \N__35503\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35547\,
            I => \N__35503\
        );

    \I__7086\ : InMux
    port map (
            O => \N__35546\,
            I => \N__35503\
        );

    \I__7085\ : InMux
    port map (
            O => \N__35545\,
            I => \N__35493\
        );

    \I__7084\ : InMux
    port map (
            O => \N__35544\,
            I => \N__35493\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35543\,
            I => \N__35493\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35542\,
            I => \N__35493\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__35537\,
            I => \N__35488\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35479\
        );

    \I__7079\ : InMux
    port map (
            O => \N__35531\,
            I => \N__35479\
        );

    \I__7078\ : InMux
    port map (
            O => \N__35528\,
            I => \N__35479\
        );

    \I__7077\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35479\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__35520\,
            I => \N__35474\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__35503\,
            I => \N__35474\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35502\,
            I => \N__35471\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__35493\,
            I => \N__35468\
        );

    \I__7072\ : InMux
    port map (
            O => \N__35492\,
            I => \N__35463\
        );

    \I__7071\ : InMux
    port map (
            O => \N__35491\,
            I => \N__35463\
        );

    \I__7070\ : Span4Mux_v
    port map (
            O => \N__35488\,
            I => \N__35460\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__35479\,
            I => \N__35455\
        );

    \I__7068\ : Span4Mux_v
    port map (
            O => \N__35474\,
            I => \N__35455\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__35471\,
            I => \N__35450\
        );

    \I__7066\ : Span4Mux_h
    port map (
            O => \N__35468\,
            I => \N__35450\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__35463\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__35460\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7063\ : Odrv4
    port map (
            O => \N__35455\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7062\ : Odrv4
    port map (
            O => \N__35450\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7061\ : InMux
    port map (
            O => \N__35441\,
            I => \N__35407\
        );

    \I__7060\ : InMux
    port map (
            O => \N__35440\,
            I => \N__35407\
        );

    \I__7059\ : InMux
    port map (
            O => \N__35439\,
            I => \N__35407\
        );

    \I__7058\ : InMux
    port map (
            O => \N__35438\,
            I => \N__35407\
        );

    \I__7057\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35407\
        );

    \I__7056\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35407\
        );

    \I__7055\ : InMux
    port map (
            O => \N__35435\,
            I => \N__35407\
        );

    \I__7054\ : InMux
    port map (
            O => \N__35434\,
            I => \N__35390\
        );

    \I__7053\ : InMux
    port map (
            O => \N__35433\,
            I => \N__35390\
        );

    \I__7052\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35390\
        );

    \I__7051\ : InMux
    port map (
            O => \N__35431\,
            I => \N__35390\
        );

    \I__7050\ : InMux
    port map (
            O => \N__35430\,
            I => \N__35390\
        );

    \I__7049\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35390\
        );

    \I__7048\ : InMux
    port map (
            O => \N__35428\,
            I => \N__35390\
        );

    \I__7047\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35390\
        );

    \I__7046\ : InMux
    port map (
            O => \N__35426\,
            I => \N__35381\
        );

    \I__7045\ : InMux
    port map (
            O => \N__35425\,
            I => \N__35381\
        );

    \I__7044\ : InMux
    port map (
            O => \N__35424\,
            I => \N__35381\
        );

    \I__7043\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35381\
        );

    \I__7042\ : CascadeMux
    port map (
            O => \N__35422\,
            I => \N__35378\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__35407\,
            I => \N__35368\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__35390\,
            I => \N__35368\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__35381\,
            I => \N__35368\
        );

    \I__7038\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35365\
        );

    \I__7037\ : InMux
    port map (
            O => \N__35377\,
            I => \N__35362\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35359\
        );

    \I__7035\ : CascadeMux
    port map (
            O => \N__35375\,
            I => \N__35356\
        );

    \I__7034\ : Span4Mux_v
    port map (
            O => \N__35368\,
            I => \N__35352\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__35365\,
            I => \N__35345\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__35362\,
            I => \N__35345\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__35359\,
            I => \N__35345\
        );

    \I__7030\ : InMux
    port map (
            O => \N__35356\,
            I => \N__35340\
        );

    \I__7029\ : InMux
    port map (
            O => \N__35355\,
            I => \N__35340\
        );

    \I__7028\ : Sp12to4
    port map (
            O => \N__35352\,
            I => \N__35335\
        );

    \I__7027\ : Span12Mux_v
    port map (
            O => \N__35345\,
            I => \N__35335\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__35340\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__7025\ : Odrv12
    port map (
            O => \N__35335\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__7024\ : CascadeMux
    port map (
            O => \N__35330\,
            I => \N__35321\
        );

    \I__7023\ : CascadeMux
    port map (
            O => \N__35329\,
            I => \N__35318\
        );

    \I__7022\ : CascadeMux
    port map (
            O => \N__35328\,
            I => \N__35315\
        );

    \I__7021\ : CascadeMux
    port map (
            O => \N__35327\,
            I => \N__35312\
        );

    \I__7020\ : CascadeMux
    port map (
            O => \N__35326\,
            I => \N__35298\
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__35325\,
            I => \N__35295\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__35324\,
            I => \N__35292\
        );

    \I__7017\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35279\
        );

    \I__7016\ : InMux
    port map (
            O => \N__35318\,
            I => \N__35279\
        );

    \I__7015\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35279\
        );

    \I__7014\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35279\
        );

    \I__7013\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35270\
        );

    \I__7012\ : InMux
    port map (
            O => \N__35310\,
            I => \N__35270\
        );

    \I__7011\ : InMux
    port map (
            O => \N__35309\,
            I => \N__35270\
        );

    \I__7010\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35270\
        );

    \I__7009\ : InMux
    port map (
            O => \N__35307\,
            I => \N__35255\
        );

    \I__7008\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35255\
        );

    \I__7007\ : InMux
    port map (
            O => \N__35305\,
            I => \N__35255\
        );

    \I__7006\ : InMux
    port map (
            O => \N__35304\,
            I => \N__35255\
        );

    \I__7005\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35255\
        );

    \I__7004\ : InMux
    port map (
            O => \N__35302\,
            I => \N__35255\
        );

    \I__7003\ : InMux
    port map (
            O => \N__35301\,
            I => \N__35255\
        );

    \I__7002\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35250\
        );

    \I__7001\ : InMux
    port map (
            O => \N__35295\,
            I => \N__35250\
        );

    \I__7000\ : InMux
    port map (
            O => \N__35292\,
            I => \N__35245\
        );

    \I__6999\ : InMux
    port map (
            O => \N__35291\,
            I => \N__35245\
        );

    \I__6998\ : InMux
    port map (
            O => \N__35290\,
            I => \N__35242\
        );

    \I__6997\ : InMux
    port map (
            O => \N__35289\,
            I => \N__35239\
        );

    \I__6996\ : InMux
    port map (
            O => \N__35288\,
            I => \N__35236\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__35279\,
            I => \N__35229\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__35270\,
            I => \N__35229\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__35255\,
            I => \N__35229\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__35250\,
            I => \N__35226\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__35245\,
            I => \N__35223\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__35242\,
            I => \N__35216\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__35239\,
            I => \N__35216\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__35236\,
            I => \N__35216\
        );

    \I__6987\ : Span4Mux_v
    port map (
            O => \N__35229\,
            I => \N__35211\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__35226\,
            I => \N__35206\
        );

    \I__6985\ : Span4Mux_h
    port map (
            O => \N__35223\,
            I => \N__35206\
        );

    \I__6984\ : Span4Mux_v
    port map (
            O => \N__35216\,
            I => \N__35203\
        );

    \I__6983\ : InMux
    port map (
            O => \N__35215\,
            I => \N__35198\
        );

    \I__6982\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35198\
        );

    \I__6981\ : Span4Mux_h
    port map (
            O => \N__35211\,
            I => \N__35195\
        );

    \I__6980\ : Span4Mux_h
    port map (
            O => \N__35206\,
            I => \N__35192\
        );

    \I__6979\ : Span4Mux_h
    port map (
            O => \N__35203\,
            I => \N__35189\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__35198\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6977\ : Odrv4
    port map (
            O => \N__35195\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__35192\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6975\ : Odrv4
    port map (
            O => \N__35189\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6974\ : CascadeMux
    port map (
            O => \N__35180\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__6973\ : CascadeMux
    port map (
            O => \N__35177\,
            I => \N__35174\
        );

    \I__6972\ : InMux
    port map (
            O => \N__35174\,
            I => \N__35171\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__35171\,
            I => \N__35166\
        );

    \I__6970\ : CascadeMux
    port map (
            O => \N__35170\,
            I => \N__35163\
        );

    \I__6969\ : InMux
    port map (
            O => \N__35169\,
            I => \N__35160\
        );

    \I__6968\ : Span4Mux_v
    port map (
            O => \N__35166\,
            I => \N__35157\
        );

    \I__6967\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35154\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__35160\,
            I => \N__35151\
        );

    \I__6965\ : Odrv4
    port map (
            O => \N__35157\,
            I => measured_delay_tr_3
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__35154\,
            I => measured_delay_tr_3
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__35151\,
            I => measured_delay_tr_3
        );

    \I__6962\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35141\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__35141\,
            I => \N__35137\
        );

    \I__6960\ : InMux
    port map (
            O => \N__35140\,
            I => \N__35134\
        );

    \I__6959\ : Span4Mux_v
    port map (
            O => \N__35137\,
            I => \N__35128\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__35134\,
            I => \N__35128\
        );

    \I__6957\ : InMux
    port map (
            O => \N__35133\,
            I => \N__35125\
        );

    \I__6956\ : Odrv4
    port map (
            O => \N__35128\,
            I => \phase_controller_inst1.stoper_tr.N_248\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__35125\,
            I => \phase_controller_inst1.stoper_tr.N_248\
        );

    \I__6954\ : CascadeMux
    port map (
            O => \N__35120\,
            I => \N__35117\
        );

    \I__6953\ : InMux
    port map (
            O => \N__35117\,
            I => \N__35114\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__35114\,
            I => \N__35110\
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__35113\,
            I => \N__35107\
        );

    \I__6950\ : Span4Mux_v
    port map (
            O => \N__35110\,
            I => \N__35104\
        );

    \I__6949\ : InMux
    port map (
            O => \N__35107\,
            I => \N__35101\
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__35104\,
            I => measured_delay_tr_1
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__35101\,
            I => measured_delay_tr_1
        );

    \I__6946\ : InMux
    port map (
            O => \N__35096\,
            I => \N__35093\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__35093\,
            I => \N__35089\
        );

    \I__6944\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35086\
        );

    \I__6943\ : Span4Mux_v
    port map (
            O => \N__35089\,
            I => \N__35082\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__35086\,
            I => \N__35079\
        );

    \I__6941\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35076\
        );

    \I__6940\ : Odrv4
    port map (
            O => \N__35082\,
            I => measured_delay_tr_11
        );

    \I__6939\ : Odrv4
    port map (
            O => \N__35079\,
            I => measured_delay_tr_11
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__35076\,
            I => measured_delay_tr_11
        );

    \I__6937\ : InMux
    port map (
            O => \N__35069\,
            I => \N__35066\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__35066\,
            I => \N__35061\
        );

    \I__6935\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35058\
        );

    \I__6934\ : InMux
    port map (
            O => \N__35064\,
            I => \N__35055\
        );

    \I__6933\ : Span4Mux_v
    port map (
            O => \N__35061\,
            I => \N__35052\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__35058\,
            I => \N__35049\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__35055\,
            I => \N__35046\
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__35052\,
            I => measured_delay_tr_9
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__35049\,
            I => measured_delay_tr_9
        );

    \I__6928\ : Odrv4
    port map (
            O => \N__35046\,
            I => measured_delay_tr_9
        );

    \I__6927\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35034\
        );

    \I__6926\ : InMux
    port map (
            O => \N__35038\,
            I => \N__35030\
        );

    \I__6925\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35027\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__35034\,
            I => \N__35024\
        );

    \I__6923\ : InMux
    port map (
            O => \N__35033\,
            I => \N__35021\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__35030\,
            I => \N__35016\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__35027\,
            I => \N__35016\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__35024\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__35021\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__6918\ : Odrv12
    port map (
            O => \N__35016\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__6917\ : InMux
    port map (
            O => \N__35009\,
            I => \N__35005\
        );

    \I__6916\ : InMux
    port map (
            O => \N__35008\,
            I => \N__35002\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__35005\,
            I => \N__34999\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__35002\,
            I => \N__34995\
        );

    \I__6913\ : Span12Mux_v
    port map (
            O => \N__34999\,
            I => \N__34992\
        );

    \I__6912\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34989\
        );

    \I__6911\ : Odrv4
    port map (
            O => \N__34995\,
            I => measured_delay_tr_6
        );

    \I__6910\ : Odrv12
    port map (
            O => \N__34992\,
            I => measured_delay_tr_6
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__34989\,
            I => measured_delay_tr_6
        );

    \I__6908\ : InMux
    port map (
            O => \N__34982\,
            I => \N__34979\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__34979\,
            I => \N__34975\
        );

    \I__6906\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34972\
        );

    \I__6905\ : Span4Mux_v
    port map (
            O => \N__34975\,
            I => \N__34966\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__34972\,
            I => \N__34966\
        );

    \I__6903\ : InMux
    port map (
            O => \N__34971\,
            I => \N__34963\
        );

    \I__6902\ : Span4Mux_v
    port map (
            O => \N__34966\,
            I => \N__34960\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__34963\,
            I => \N__34957\
        );

    \I__6900\ : Odrv4
    port map (
            O => \N__34960\,
            I => measured_delay_tr_2
        );

    \I__6899\ : Odrv4
    port map (
            O => \N__34957\,
            I => measured_delay_tr_2
        );

    \I__6898\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34948\
        );

    \I__6897\ : InMux
    port map (
            O => \N__34951\,
            I => \N__34945\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__34948\,
            I => \N__34940\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34945\,
            I => \N__34940\
        );

    \I__6894\ : Span4Mux_v
    port map (
            O => \N__34940\,
            I => \N__34935\
        );

    \I__6893\ : InMux
    port map (
            O => \N__34939\,
            I => \N__34932\
        );

    \I__6892\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34929\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__34935\,
            I => \phase_controller_inst1.stoper_tr.N_55\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__34932\,
            I => \phase_controller_inst1.stoper_tr.N_55\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__34929\,
            I => \phase_controller_inst1.stoper_tr.N_55\
        );

    \I__6888\ : InMux
    port map (
            O => \N__34922\,
            I => \N__34919\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__34919\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\
        );

    \I__6886\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34913\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__34913\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\
        );

    \I__6884\ : InMux
    port map (
            O => \N__34910\,
            I => \N__34907\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__34907\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\
        );

    \I__6882\ : CascadeMux
    port map (
            O => \N__34904\,
            I => \N__34901\
        );

    \I__6881\ : InMux
    port map (
            O => \N__34901\,
            I => \N__34898\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__34898\,
            I => \N__34895\
        );

    \I__6879\ : Odrv12
    port map (
            O => \N__34895\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__6878\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34889\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__34889\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\
        );

    \I__6876\ : InMux
    port map (
            O => \N__34886\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__6875\ : CascadeMux
    port map (
            O => \N__34883\,
            I => \N__34880\
        );

    \I__6874\ : InMux
    port map (
            O => \N__34880\,
            I => \N__34877\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__34877\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__6872\ : CascadeMux
    port map (
            O => \N__34874\,
            I => \N__34871\
        );

    \I__6871\ : InMux
    port map (
            O => \N__34871\,
            I => \N__34868\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__34868\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__6869\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34861\
        );

    \I__6868\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34857\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__34861\,
            I => \N__34854\
        );

    \I__6866\ : InMux
    port map (
            O => \N__34860\,
            I => \N__34851\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__34857\,
            I => \N__34848\
        );

    \I__6864\ : Odrv4
    port map (
            O => \N__34854\,
            I => measured_delay_tr_5
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__34851\,
            I => measured_delay_tr_5
        );

    \I__6862\ : Odrv4
    port map (
            O => \N__34848\,
            I => measured_delay_tr_5
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__34841\,
            I => \N__34838\
        );

    \I__6860\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34835\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__34835\,
            I => \N__34832\
        );

    \I__6858\ : Odrv12
    port map (
            O => \N__34832\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__6857\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34826\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__34826\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__6855\ : CascadeMux
    port map (
            O => \N__34823\,
            I => \N__34820\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34817\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__34817\,
            I => \N__34814\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__34814\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__6851\ : InMux
    port map (
            O => \N__34811\,
            I => \N__34808\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__34808\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__6849\ : InMux
    port map (
            O => \N__34805\,
            I => \N__34802\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__34802\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__6847\ : CascadeMux
    port map (
            O => \N__34799\,
            I => \N__34796\
        );

    \I__6846\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34793\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__34793\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34790\,
            I => \N__34787\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34787\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__6842\ : CascadeMux
    port map (
            O => \N__34784\,
            I => \N__34781\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34781\,
            I => \N__34778\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__34778\,
            I => \N__34775\
        );

    \I__6839\ : Span4Mux_h
    port map (
            O => \N__34775\,
            I => \N__34772\
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__34772\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__6837\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34766\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__34766\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__6835\ : InMux
    port map (
            O => \N__34763\,
            I => \N__34760\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34760\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__6833\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34754\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__34754\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__6831\ : CascadeMux
    port map (
            O => \N__34751\,
            I => \N__34748\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34748\,
            I => \N__34745\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__34745\,
            I => \N__34742\
        );

    \I__6828\ : Span4Mux_v
    port map (
            O => \N__34742\,
            I => \N__34739\
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__34739\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__6826\ : InMux
    port map (
            O => \N__34736\,
            I => \N__34733\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__34733\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__6824\ : InMux
    port map (
            O => \N__34730\,
            I => \N__34727\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__34727\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__6822\ : CascadeMux
    port map (
            O => \N__34724\,
            I => \N__34721\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34721\,
            I => \N__34718\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__34718\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__6819\ : CascadeMux
    port map (
            O => \N__34715\,
            I => \N__34712\
        );

    \I__6818\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34709\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__34709\,
            I => \N__34706\
        );

    \I__6816\ : Odrv4
    port map (
            O => \N__34706\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__6815\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34700\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__34700\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__34697\,
            I => \N__34694\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34691\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__34691\,
            I => \N__34688\
        );

    \I__6810\ : Odrv12
    port map (
            O => \N__34688\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34682\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__34682\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34676\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__34676\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__6805\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34670\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__34670\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__34667\,
            I => \N__34664\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34664\,
            I => \N__34661\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__34661\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__6800\ : CascadeMux
    port map (
            O => \N__34658\,
            I => \N__34655\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34652\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__34652\,
            I => \N__34649\
        );

    \I__6797\ : Span4Mux_h
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__34646\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__6795\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34640\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34640\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__34637\,
            I => \N__34634\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34631\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34631\,
            I => \N__34628\
        );

    \I__6790\ : Span4Mux_h
    port map (
            O => \N__34628\,
            I => \N__34625\
        );

    \I__6789\ : Odrv4
    port map (
            O => \N__34625\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34622\,
            I => \N__34619\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34619\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__6786\ : CascadeMux
    port map (
            O => \N__34616\,
            I => \N__34613\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34603\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34603\
        );

    \I__6783\ : CascadeMux
    port map (
            O => \N__34611\,
            I => \N__34600\
        );

    \I__6782\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34593\
        );

    \I__6781\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34593\
        );

    \I__6780\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34593\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__34603\,
            I => \N__34590\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34587\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__34593\,
            I => \N__34584\
        );

    \I__6776\ : Span4Mux_h
    port map (
            O => \N__34590\,
            I => \N__34581\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__34587\,
            I => state_3
        );

    \I__6774\ : Odrv12
    port map (
            O => \N__34584\,
            I => state_3
        );

    \I__6773\ : Odrv4
    port map (
            O => \N__34581\,
            I => state_3
        );

    \I__6772\ : IoInMux
    port map (
            O => \N__34574\,
            I => \N__34571\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__34571\,
            I => \N__34568\
        );

    \I__6770\ : Span4Mux_s1_v
    port map (
            O => \N__34568\,
            I => \N__34564\
        );

    \I__6769\ : CascadeMux
    port map (
            O => \N__34567\,
            I => \N__34561\
        );

    \I__6768\ : Span4Mux_v
    port map (
            O => \N__34564\,
            I => \N__34557\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34552\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34552\
        );

    \I__6765\ : Odrv4
    port map (
            O => \N__34557\,
            I => s1_phy_c
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__34552\,
            I => s1_phy_c
        );

    \I__6763\ : InMux
    port map (
            O => \N__34547\,
            I => \N__34537\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34546\,
            I => \N__34537\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34545\,
            I => \N__34537\
        );

    \I__6760\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34534\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__34537\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__34534\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6757\ : IoInMux
    port map (
            O => \N__34529\,
            I => \N__34526\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__34526\,
            I => \N__34523\
        );

    \I__6755\ : Odrv12
    port map (
            O => \N__34523\,
            I => \current_shift_inst.timer_s1.N_181_i\
        );

    \I__6754\ : IoInMux
    port map (
            O => \N__34520\,
            I => \N__34517\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__34517\,
            I => \N__34514\
        );

    \I__6752\ : Odrv12
    port map (
            O => \N__34514\,
            I => s2_phy_c
        );

    \I__6751\ : CascadeMux
    port map (
            O => \N__34511\,
            I => \phase_controller_inst2.stoper_tr.time_passed11_cascade_\
        );

    \I__6750\ : CascadeMux
    port map (
            O => \N__34508\,
            I => \N__34503\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34507\,
            I => \N__34499\
        );

    \I__6748\ : CascadeMux
    port map (
            O => \N__34506\,
            I => \N__34496\
        );

    \I__6747\ : InMux
    port map (
            O => \N__34503\,
            I => \N__34493\
        );

    \I__6746\ : CascadeMux
    port map (
            O => \N__34502\,
            I => \N__34490\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__34499\,
            I => \N__34487\
        );

    \I__6744\ : InMux
    port map (
            O => \N__34496\,
            I => \N__34484\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__34493\,
            I => \N__34481\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34478\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__34487\,
            I => \N__34475\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__34484\,
            I => \N__34472\
        );

    \I__6739\ : Span4Mux_h
    port map (
            O => \N__34481\,
            I => \N__34467\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__34478\,
            I => \N__34467\
        );

    \I__6737\ : Span4Mux_v
    port map (
            O => \N__34475\,
            I => \N__34463\
        );

    \I__6736\ : Span4Mux_h
    port map (
            O => \N__34472\,
            I => \N__34458\
        );

    \I__6735\ : Span4Mux_h
    port map (
            O => \N__34467\,
            I => \N__34458\
        );

    \I__6734\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34455\
        );

    \I__6733\ : Span4Mux_h
    port map (
            O => \N__34463\,
            I => \N__34452\
        );

    \I__6732\ : Span4Mux_v
    port map (
            O => \N__34458\,
            I => \N__34449\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__34455\,
            I => measured_delay_hc_13
        );

    \I__6730\ : Odrv4
    port map (
            O => \N__34452\,
            I => measured_delay_hc_13
        );

    \I__6729\ : Odrv4
    port map (
            O => \N__34449\,
            I => measured_delay_hc_13
        );

    \I__6728\ : CascadeMux
    port map (
            O => \N__34442\,
            I => \N__34439\
        );

    \I__6727\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34436\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__34436\,
            I => \N__34433\
        );

    \I__6725\ : Odrv12
    port map (
            O => \N__34433\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34425\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34421\
        );

    \I__6722\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34418\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__34425\,
            I => \N__34415\
        );

    \I__6720\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34412\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__34421\,
            I => \N__34409\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__34418\,
            I => \N__34406\
        );

    \I__6717\ : Span4Mux_h
    port map (
            O => \N__34415\,
            I => \N__34401\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__34412\,
            I => \N__34401\
        );

    \I__6715\ : Span4Mux_h
    port map (
            O => \N__34409\,
            I => \N__34395\
        );

    \I__6714\ : Span4Mux_h
    port map (
            O => \N__34406\,
            I => \N__34395\
        );

    \I__6713\ : Span4Mux_h
    port map (
            O => \N__34401\,
            I => \N__34392\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34400\,
            I => \N__34389\
        );

    \I__6711\ : Span4Mux_v
    port map (
            O => \N__34395\,
            I => \N__34386\
        );

    \I__6710\ : Odrv4
    port map (
            O => \N__34392\,
            I => measured_delay_hc_15
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__34389\,
            I => measured_delay_hc_15
        );

    \I__6708\ : Odrv4
    port map (
            O => \N__34386\,
            I => measured_delay_hc_15
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__34379\,
            I => \N__34376\
        );

    \I__6706\ : InMux
    port map (
            O => \N__34376\,
            I => \N__34373\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__34373\,
            I => \N__34370\
        );

    \I__6704\ : Span4Mux_v
    port map (
            O => \N__34370\,
            I => \N__34367\
        );

    \I__6703\ : Odrv4
    port map (
            O => \N__34367\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__6702\ : CascadeMux
    port map (
            O => \N__34364\,
            I => \N__34353\
        );

    \I__6701\ : CascadeMux
    port map (
            O => \N__34363\,
            I => \N__34350\
        );

    \I__6700\ : CascadeMux
    port map (
            O => \N__34362\,
            I => \N__34347\
        );

    \I__6699\ : CascadeMux
    port map (
            O => \N__34361\,
            I => \N__34344\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34360\,
            I => \N__34329\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34359\,
            I => \N__34329\
        );

    \I__6696\ : InMux
    port map (
            O => \N__34358\,
            I => \N__34329\
        );

    \I__6695\ : InMux
    port map (
            O => \N__34357\,
            I => \N__34326\
        );

    \I__6694\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34309\
        );

    \I__6693\ : InMux
    port map (
            O => \N__34353\,
            I => \N__34309\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34350\,
            I => \N__34309\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34309\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34344\,
            I => \N__34309\
        );

    \I__6689\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34309\
        );

    \I__6688\ : InMux
    port map (
            O => \N__34342\,
            I => \N__34309\
        );

    \I__6687\ : InMux
    port map (
            O => \N__34341\,
            I => \N__34309\
        );

    \I__6686\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34304\
        );

    \I__6685\ : InMux
    port map (
            O => \N__34339\,
            I => \N__34304\
        );

    \I__6684\ : CascadeMux
    port map (
            O => \N__34338\,
            I => \N__34300\
        );

    \I__6683\ : CascadeMux
    port map (
            O => \N__34337\,
            I => \N__34297\
        );

    \I__6682\ : CascadeMux
    port map (
            O => \N__34336\,
            I => \N__34285\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__34329\,
            I => \N__34277\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__34326\,
            I => \N__34277\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__34309\,
            I => \N__34277\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__34304\,
            I => \N__34274\
        );

    \I__6677\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34271\
        );

    \I__6676\ : InMux
    port map (
            O => \N__34300\,
            I => \N__34259\
        );

    \I__6675\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34259\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34250\
        );

    \I__6673\ : InMux
    port map (
            O => \N__34295\,
            I => \N__34250\
        );

    \I__6672\ : InMux
    port map (
            O => \N__34294\,
            I => \N__34250\
        );

    \I__6671\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34250\
        );

    \I__6670\ : InMux
    port map (
            O => \N__34292\,
            I => \N__34239\
        );

    \I__6669\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34239\
        );

    \I__6668\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34239\
        );

    \I__6667\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34239\
        );

    \I__6666\ : InMux
    port map (
            O => \N__34288\,
            I => \N__34239\
        );

    \I__6665\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34234\
        );

    \I__6664\ : InMux
    port map (
            O => \N__34284\,
            I => \N__34234\
        );

    \I__6663\ : Span4Mux_v
    port map (
            O => \N__34277\,
            I => \N__34227\
        );

    \I__6662\ : Span4Mux_v
    port map (
            O => \N__34274\,
            I => \N__34227\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__34271\,
            I => \N__34227\
        );

    \I__6660\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34224\
        );

    \I__6659\ : InMux
    port map (
            O => \N__34269\,
            I => \N__34211\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34268\,
            I => \N__34211\
        );

    \I__6657\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34211\
        );

    \I__6656\ : InMux
    port map (
            O => \N__34266\,
            I => \N__34211\
        );

    \I__6655\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34211\
        );

    \I__6654\ : InMux
    port map (
            O => \N__34264\,
            I => \N__34211\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__34259\,
            I => \N__34206\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__34250\,
            I => \N__34206\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__34239\,
            I => \N__34203\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__34234\,
            I => \N__34200\
        );

    \I__6649\ : Span4Mux_h
    port map (
            O => \N__34227\,
            I => \N__34197\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__34224\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__34211\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\
        );

    \I__6646\ : Odrv4
    port map (
            O => \N__34206\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\
        );

    \I__6645\ : Odrv4
    port map (
            O => \N__34203\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\
        );

    \I__6644\ : Odrv12
    port map (
            O => \N__34200\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\
        );

    \I__6643\ : Odrv4
    port map (
            O => \N__34197\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\
        );

    \I__6642\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34178\
        );

    \I__6641\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34178\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__34178\,
            I => \N__34162\
        );

    \I__6639\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34157\
        );

    \I__6638\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34157\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34175\,
            I => \N__34142\
        );

    \I__6636\ : InMux
    port map (
            O => \N__34174\,
            I => \N__34142\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34142\
        );

    \I__6634\ : InMux
    port map (
            O => \N__34172\,
            I => \N__34142\
        );

    \I__6633\ : InMux
    port map (
            O => \N__34171\,
            I => \N__34142\
        );

    \I__6632\ : InMux
    port map (
            O => \N__34170\,
            I => \N__34142\
        );

    \I__6631\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34131\
        );

    \I__6630\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34131\
        );

    \I__6629\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34131\
        );

    \I__6628\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34131\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34131\
        );

    \I__6626\ : Span4Mux_h
    port map (
            O => \N__34162\,
            I => \N__34123\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__34157\,
            I => \N__34123\
        );

    \I__6624\ : InMux
    port map (
            O => \N__34156\,
            I => \N__34118\
        );

    \I__6623\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34118\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__34142\,
            I => \N__34115\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__34131\,
            I => \N__34112\
        );

    \I__6620\ : InMux
    port map (
            O => \N__34130\,
            I => \N__34105\
        );

    \I__6619\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34105\
        );

    \I__6618\ : InMux
    port map (
            O => \N__34128\,
            I => \N__34105\
        );

    \I__6617\ : Span4Mux_h
    port map (
            O => \N__34123\,
            I => \N__34094\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__34118\,
            I => \N__34091\
        );

    \I__6615\ : Span4Mux_v
    port map (
            O => \N__34115\,
            I => \N__34084\
        );

    \I__6614\ : Span4Mux_h
    port map (
            O => \N__34112\,
            I => \N__34084\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__34105\,
            I => \N__34084\
        );

    \I__6612\ : InMux
    port map (
            O => \N__34104\,
            I => \N__34067\
        );

    \I__6611\ : InMux
    port map (
            O => \N__34103\,
            I => \N__34067\
        );

    \I__6610\ : InMux
    port map (
            O => \N__34102\,
            I => \N__34067\
        );

    \I__6609\ : InMux
    port map (
            O => \N__34101\,
            I => \N__34067\
        );

    \I__6608\ : InMux
    port map (
            O => \N__34100\,
            I => \N__34067\
        );

    \I__6607\ : InMux
    port map (
            O => \N__34099\,
            I => \N__34067\
        );

    \I__6606\ : InMux
    port map (
            O => \N__34098\,
            I => \N__34067\
        );

    \I__6605\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34067\
        );

    \I__6604\ : Odrv4
    port map (
            O => \N__34094\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt30\
        );

    \I__6603\ : Odrv4
    port map (
            O => \N__34091\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt30\
        );

    \I__6602\ : Odrv4
    port map (
            O => \N__34084\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt30\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__34067\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt30\
        );

    \I__6600\ : CascadeMux
    port map (
            O => \N__34058\,
            I => \N__34055\
        );

    \I__6599\ : InMux
    port map (
            O => \N__34055\,
            I => \N__34051\
        );

    \I__6598\ : CascadeMux
    port map (
            O => \N__34054\,
            I => \N__34048\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__34051\,
            I => \N__34045\
        );

    \I__6596\ : InMux
    port map (
            O => \N__34048\,
            I => \N__34040\
        );

    \I__6595\ : Span4Mux_v
    port map (
            O => \N__34045\,
            I => \N__34036\
        );

    \I__6594\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34031\
        );

    \I__6593\ : InMux
    port map (
            O => \N__34043\,
            I => \N__34031\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__34040\,
            I => \N__34028\
        );

    \I__6591\ : InMux
    port map (
            O => \N__34039\,
            I => \N__34025\
        );

    \I__6590\ : Span4Mux_h
    port map (
            O => \N__34036\,
            I => \N__34020\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__34031\,
            I => \N__34020\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__34028\,
            I => measured_delay_hc_2
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__34025\,
            I => measured_delay_hc_2
        );

    \I__6586\ : Odrv4
    port map (
            O => \N__34020\,
            I => measured_delay_hc_2
        );

    \I__6585\ : CascadeMux
    port map (
            O => \N__34013\,
            I => \N__34005\
        );

    \I__6584\ : CascadeMux
    port map (
            O => \N__34012\,
            I => \N__33999\
        );

    \I__6583\ : CascadeMux
    port map (
            O => \N__34011\,
            I => \N__33996\
        );

    \I__6582\ : CascadeMux
    port map (
            O => \N__34010\,
            I => \N__33993\
        );

    \I__6581\ : InMux
    port map (
            O => \N__34009\,
            I => \N__33987\
        );

    \I__6580\ : InMux
    port map (
            O => \N__34008\,
            I => \N__33987\
        );

    \I__6579\ : InMux
    port map (
            O => \N__34005\,
            I => \N__33976\
        );

    \I__6578\ : InMux
    port map (
            O => \N__34004\,
            I => \N__33976\
        );

    \I__6577\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33976\
        );

    \I__6576\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33976\
        );

    \I__6575\ : InMux
    port map (
            O => \N__33999\,
            I => \N__33967\
        );

    \I__6574\ : InMux
    port map (
            O => \N__33996\,
            I => \N__33967\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33993\,
            I => \N__33967\
        );

    \I__6572\ : InMux
    port map (
            O => \N__33992\,
            I => \N__33967\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__33987\,
            I => \N__33964\
        );

    \I__6570\ : CascadeMux
    port map (
            O => \N__33986\,
            I => \N__33952\
        );

    \I__6569\ : CascadeMux
    port map (
            O => \N__33985\,
            I => \N__33949\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__33976\,
            I => \N__33942\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__33967\,
            I => \N__33937\
        );

    \I__6566\ : Span4Mux_h
    port map (
            O => \N__33964\,
            I => \N__33937\
        );

    \I__6565\ : CascadeMux
    port map (
            O => \N__33963\,
            I => \N__33932\
        );

    \I__6564\ : CascadeMux
    port map (
            O => \N__33962\,
            I => \N__33929\
        );

    \I__6563\ : CascadeMux
    port map (
            O => \N__33961\,
            I => \N__33924\
        );

    \I__6562\ : CascadeMux
    port map (
            O => \N__33960\,
            I => \N__33918\
        );

    \I__6561\ : CascadeMux
    port map (
            O => \N__33959\,
            I => \N__33915\
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__33958\,
            I => \N__33912\
        );

    \I__6559\ : InMux
    port map (
            O => \N__33957\,
            I => \N__33904\
        );

    \I__6558\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33887\
        );

    \I__6557\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33887\
        );

    \I__6556\ : InMux
    port map (
            O => \N__33952\,
            I => \N__33887\
        );

    \I__6555\ : InMux
    port map (
            O => \N__33949\,
            I => \N__33887\
        );

    \I__6554\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33887\
        );

    \I__6553\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33887\
        );

    \I__6552\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33887\
        );

    \I__6551\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33887\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__33942\,
            I => \N__33884\
        );

    \I__6549\ : Span4Mux_h
    port map (
            O => \N__33937\,
            I => \N__33881\
        );

    \I__6548\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33878\
        );

    \I__6547\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33867\
        );

    \I__6546\ : InMux
    port map (
            O => \N__33932\,
            I => \N__33867\
        );

    \I__6545\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33867\
        );

    \I__6544\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33867\
        );

    \I__6543\ : InMux
    port map (
            O => \N__33927\,
            I => \N__33867\
        );

    \I__6542\ : InMux
    port map (
            O => \N__33924\,
            I => \N__33858\
        );

    \I__6541\ : InMux
    port map (
            O => \N__33923\,
            I => \N__33858\
        );

    \I__6540\ : InMux
    port map (
            O => \N__33922\,
            I => \N__33858\
        );

    \I__6539\ : InMux
    port map (
            O => \N__33921\,
            I => \N__33858\
        );

    \I__6538\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33841\
        );

    \I__6537\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33841\
        );

    \I__6536\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33841\
        );

    \I__6535\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33841\
        );

    \I__6534\ : InMux
    port map (
            O => \N__33910\,
            I => \N__33841\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33909\,
            I => \N__33841\
        );

    \I__6532\ : InMux
    port map (
            O => \N__33908\,
            I => \N__33841\
        );

    \I__6531\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33841\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__33904\,
            I => \N__33836\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__33887\,
            I => \N__33836\
        );

    \I__6528\ : Span4Mux_h
    port map (
            O => \N__33884\,
            I => \N__33831\
        );

    \I__6527\ : Span4Mux_h
    port map (
            O => \N__33881\,
            I => \N__33831\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__33878\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__33867\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__33858\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__33841\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6522\ : Odrv12
    port map (
            O => \N__33836\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6521\ : Odrv4
    port map (
            O => \N__33831\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6520\ : CascadeMux
    port map (
            O => \N__33818\,
            I => \N__33815\
        );

    \I__6519\ : InMux
    port map (
            O => \N__33815\,
            I => \N__33812\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__33812\,
            I => \N__33809\
        );

    \I__6517\ : Span4Mux_v
    port map (
            O => \N__33809\,
            I => \N__33806\
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__33806\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__6515\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33800\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__33800\,
            I => \N__33795\
        );

    \I__6513\ : InMux
    port map (
            O => \N__33799\,
            I => \N__33790\
        );

    \I__6512\ : InMux
    port map (
            O => \N__33798\,
            I => \N__33790\
        );

    \I__6511\ : Span12Mux_h
    port map (
            O => \N__33795\,
            I => \N__33787\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__33790\,
            I => \N__33784\
        );

    \I__6509\ : Span12Mux_v
    port map (
            O => \N__33787\,
            I => \N__33781\
        );

    \I__6508\ : Span12Mux_v
    port map (
            O => \N__33784\,
            I => \N__33778\
        );

    \I__6507\ : Odrv12
    port map (
            O => \N__33781\,
            I => \il_max_comp1_D2\
        );

    \I__6506\ : Odrv12
    port map (
            O => \N__33778\,
            I => \il_max_comp1_D2\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33773\,
            I => \N__33770\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__33770\,
            I => \N__33766\
        );

    \I__6503\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33763\
        );

    \I__6502\ : Span4Mux_h
    port map (
            O => \N__33766\,
            I => \N__33758\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__33763\,
            I => \N__33758\
        );

    \I__6500\ : Odrv4
    port map (
            O => \N__33758\,
            I => state_ns_i_a3_1
        );

    \I__6499\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33752\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__33752\,
            I => \N__33747\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33751\,
            I => \N__33744\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33740\
        );

    \I__6495\ : Span4Mux_v
    port map (
            O => \N__33747\,
            I => \N__33735\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__33744\,
            I => \N__33735\
        );

    \I__6493\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33732\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__33740\,
            I => \N__33729\
        );

    \I__6491\ : Span4Mux_v
    port map (
            O => \N__33735\,
            I => \N__33725\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__33732\,
            I => \N__33720\
        );

    \I__6489\ : Span4Mux_h
    port map (
            O => \N__33729\,
            I => \N__33720\
        );

    \I__6488\ : InMux
    port map (
            O => \N__33728\,
            I => \N__33717\
        );

    \I__6487\ : Span4Mux_h
    port map (
            O => \N__33725\,
            I => \N__33714\
        );

    \I__6486\ : Span4Mux_v
    port map (
            O => \N__33720\,
            I => \N__33711\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__33717\,
            I => measured_delay_hc_12
        );

    \I__6484\ : Odrv4
    port map (
            O => \N__33714\,
            I => measured_delay_hc_12
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__33711\,
            I => measured_delay_hc_12
        );

    \I__6482\ : InMux
    port map (
            O => \N__33704\,
            I => \N__33699\
        );

    \I__6481\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33695\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33702\,
            I => \N__33692\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__33699\,
            I => \N__33689\
        );

    \I__6478\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33686\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__33695\,
            I => \N__33682\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__33692\,
            I => \N__33679\
        );

    \I__6475\ : Span4Mux_h
    port map (
            O => \N__33689\,
            I => \N__33674\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__33686\,
            I => \N__33674\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33685\,
            I => \N__33671\
        );

    \I__6472\ : Span4Mux_h
    port map (
            O => \N__33682\,
            I => \N__33668\
        );

    \I__6471\ : Span4Mux_v
    port map (
            O => \N__33679\,
            I => \N__33665\
        );

    \I__6470\ : Span4Mux_h
    port map (
            O => \N__33674\,
            I => \N__33662\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__33671\,
            I => \N__33659\
        );

    \I__6468\ : Span4Mux_v
    port map (
            O => \N__33668\,
            I => \N__33654\
        );

    \I__6467\ : Span4Mux_h
    port map (
            O => \N__33665\,
            I => \N__33654\
        );

    \I__6466\ : Span4Mux_v
    port map (
            O => \N__33662\,
            I => \N__33651\
        );

    \I__6465\ : Odrv4
    port map (
            O => \N__33659\,
            I => measured_delay_hc_11
        );

    \I__6464\ : Odrv4
    port map (
            O => \N__33654\,
            I => measured_delay_hc_11
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__33651\,
            I => measured_delay_hc_11
        );

    \I__6462\ : CascadeMux
    port map (
            O => \N__33644\,
            I => \N__33639\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33636\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__33642\,
            I => \N__33632\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33639\,
            I => \N__33629\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__33636\,
            I => \N__33626\
        );

    \I__6457\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33623\
        );

    \I__6456\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33620\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__33629\,
            I => \N__33616\
        );

    \I__6454\ : Span4Mux_v
    port map (
            O => \N__33626\,
            I => \N__33611\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__33623\,
            I => \N__33611\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__33620\,
            I => \N__33608\
        );

    \I__6451\ : InMux
    port map (
            O => \N__33619\,
            I => \N__33605\
        );

    \I__6450\ : Span4Mux_v
    port map (
            O => \N__33616\,
            I => \N__33598\
        );

    \I__6449\ : Span4Mux_v
    port map (
            O => \N__33611\,
            I => \N__33598\
        );

    \I__6448\ : Span4Mux_v
    port map (
            O => \N__33608\,
            I => \N__33598\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__33605\,
            I => measured_delay_hc_9
        );

    \I__6446\ : Odrv4
    port map (
            O => \N__33598\,
            I => measured_delay_hc_9
        );

    \I__6445\ : CascadeMux
    port map (
            O => \N__33593\,
            I => \N__33589\
        );

    \I__6444\ : CascadeMux
    port map (
            O => \N__33592\,
            I => \N__33586\
        );

    \I__6443\ : InMux
    port map (
            O => \N__33589\,
            I => \N__33582\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33578\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33575\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__33582\,
            I => \N__33571\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33568\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__33578\,
            I => \N__33565\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33575\,
            I => \N__33562\
        );

    \I__6436\ : InMux
    port map (
            O => \N__33574\,
            I => \N__33559\
        );

    \I__6435\ : Span4Mux_v
    port map (
            O => \N__33571\,
            I => \N__33556\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__33568\,
            I => \N__33553\
        );

    \I__6433\ : Span4Mux_v
    port map (
            O => \N__33565\,
            I => \N__33548\
        );

    \I__6432\ : Span4Mux_v
    port map (
            O => \N__33562\,
            I => \N__33548\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__33559\,
            I => \N__33545\
        );

    \I__6430\ : Span4Mux_h
    port map (
            O => \N__33556\,
            I => \N__33540\
        );

    \I__6429\ : Span4Mux_v
    port map (
            O => \N__33553\,
            I => \N__33540\
        );

    \I__6428\ : Odrv4
    port map (
            O => \N__33548\,
            I => measured_delay_hc_10
        );

    \I__6427\ : Odrv12
    port map (
            O => \N__33545\,
            I => measured_delay_hc_10
        );

    \I__6426\ : Odrv4
    port map (
            O => \N__33540\,
            I => measured_delay_hc_10
        );

    \I__6425\ : InMux
    port map (
            O => \N__33533\,
            I => \N__33530\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33530\,
            I => \N__33527\
        );

    \I__6423\ : Odrv4
    port map (
            O => \N__33527\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\
        );

    \I__6422\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33504\
        );

    \I__6421\ : CascadeMux
    port map (
            O => \N__33523\,
            I => \N__33501\
        );

    \I__6420\ : CascadeMux
    port map (
            O => \N__33522\,
            I => \N__33496\
        );

    \I__6419\ : InMux
    port map (
            O => \N__33521\,
            I => \N__33491\
        );

    \I__6418\ : InMux
    port map (
            O => \N__33520\,
            I => \N__33491\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33519\,
            I => \N__33482\
        );

    \I__6416\ : InMux
    port map (
            O => \N__33518\,
            I => \N__33482\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33517\,
            I => \N__33482\
        );

    \I__6414\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33482\
        );

    \I__6413\ : InMux
    port map (
            O => \N__33515\,
            I => \N__33479\
        );

    \I__6412\ : InMux
    port map (
            O => \N__33514\,
            I => \N__33470\
        );

    \I__6411\ : InMux
    port map (
            O => \N__33513\,
            I => \N__33465\
        );

    \I__6410\ : InMux
    port map (
            O => \N__33512\,
            I => \N__33465\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33511\,
            I => \N__33460\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33460\
        );

    \I__6407\ : InMux
    port map (
            O => \N__33509\,
            I => \N__33453\
        );

    \I__6406\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33453\
        );

    \I__6405\ : InMux
    port map (
            O => \N__33507\,
            I => \N__33453\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__33504\,
            I => \N__33448\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33443\
        );

    \I__6402\ : InMux
    port map (
            O => \N__33500\,
            I => \N__33443\
        );

    \I__6401\ : InMux
    port map (
            O => \N__33499\,
            I => \N__33438\
        );

    \I__6400\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33438\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__33491\,
            I => \N__33432\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__33482\,
            I => \N__33432\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__33479\,
            I => \N__33429\
        );

    \I__6396\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33418\
        );

    \I__6395\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33418\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33418\
        );

    \I__6393\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33418\
        );

    \I__6392\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33418\
        );

    \I__6391\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33415\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__33470\,
            I => \N__33411\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__33465\,
            I => \N__33408\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__33460\,
            I => \N__33405\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__33453\,
            I => \N__33402\
        );

    \I__6386\ : InMux
    port map (
            O => \N__33452\,
            I => \N__33397\
        );

    \I__6385\ : InMux
    port map (
            O => \N__33451\,
            I => \N__33397\
        );

    \I__6384\ : Span4Mux_v
    port map (
            O => \N__33448\,
            I => \N__33392\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__33443\,
            I => \N__33392\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__33438\,
            I => \N__33389\
        );

    \I__6381\ : InMux
    port map (
            O => \N__33437\,
            I => \N__33386\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__33432\,
            I => \N__33379\
        );

    \I__6379\ : Span4Mux_h
    port map (
            O => \N__33429\,
            I => \N__33379\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__33418\,
            I => \N__33379\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__33415\,
            I => \N__33373\
        );

    \I__6376\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33370\
        );

    \I__6375\ : Span4Mux_v
    port map (
            O => \N__33411\,
            I => \N__33359\
        );

    \I__6374\ : Span4Mux_v
    port map (
            O => \N__33408\,
            I => \N__33359\
        );

    \I__6373\ : Span4Mux_v
    port map (
            O => \N__33405\,
            I => \N__33359\
        );

    \I__6372\ : Span4Mux_v
    port map (
            O => \N__33402\,
            I => \N__33359\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__33397\,
            I => \N__33359\
        );

    \I__6370\ : Span4Mux_h
    port map (
            O => \N__33392\,
            I => \N__33354\
        );

    \I__6369\ : Span4Mux_h
    port map (
            O => \N__33389\,
            I => \N__33354\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__33386\,
            I => \N__33349\
        );

    \I__6367\ : Span4Mux_h
    port map (
            O => \N__33379\,
            I => \N__33349\
        );

    \I__6366\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33344\
        );

    \I__6365\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33344\
        );

    \I__6364\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33341\
        );

    \I__6363\ : Odrv4
    port map (
            O => \N__33373\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__33370\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__6361\ : Odrv4
    port map (
            O => \N__33359\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__6360\ : Odrv4
    port map (
            O => \N__33354\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__33349\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__33344\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__33341\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__6356\ : CascadeMux
    port map (
            O => \N__33326\,
            I => \N__33309\
        );

    \I__6355\ : InMux
    port map (
            O => \N__33325\,
            I => \N__33302\
        );

    \I__6354\ : InMux
    port map (
            O => \N__33324\,
            I => \N__33302\
        );

    \I__6353\ : InMux
    port map (
            O => \N__33323\,
            I => \N__33297\
        );

    \I__6352\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33297\
        );

    \I__6351\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33294\
        );

    \I__6350\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33290\
        );

    \I__6349\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33286\
        );

    \I__6348\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33283\
        );

    \I__6347\ : InMux
    port map (
            O => \N__33317\,
            I => \N__33280\
        );

    \I__6346\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33277\
        );

    \I__6345\ : InMux
    port map (
            O => \N__33315\,
            I => \N__33274\
        );

    \I__6344\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33268\
        );

    \I__6343\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33263\
        );

    \I__6342\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33263\
        );

    \I__6341\ : InMux
    port map (
            O => \N__33309\,
            I => \N__33252\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33308\,
            I => \N__33252\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33252\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__33302\,
            I => \N__33245\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__33297\,
            I => \N__33245\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__33294\,
            I => \N__33245\
        );

    \I__6335\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33242\
        );

    \I__6334\ : LocalMux
    port map (
            O => \N__33290\,
            I => \N__33239\
        );

    \I__6333\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33236\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__33286\,
            I => \N__33231\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__33283\,
            I => \N__33231\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__33280\,
            I => \N__33224\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__33277\,
            I => \N__33224\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__33274\,
            I => \N__33224\
        );

    \I__6327\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33217\
        );

    \I__6326\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33217\
        );

    \I__6325\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33217\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__33268\,
            I => \N__33212\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__33263\,
            I => \N__33212\
        );

    \I__6322\ : InMux
    port map (
            O => \N__33262\,
            I => \N__33207\
        );

    \I__6321\ : InMux
    port map (
            O => \N__33261\,
            I => \N__33207\
        );

    \I__6320\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33197\
        );

    \I__6319\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33197\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__33252\,
            I => \N__33188\
        );

    \I__6317\ : Span4Mux_v
    port map (
            O => \N__33245\,
            I => \N__33188\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__33242\,
            I => \N__33188\
        );

    \I__6315\ : Span4Mux_v
    port map (
            O => \N__33239\,
            I => \N__33188\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__33236\,
            I => \N__33185\
        );

    \I__6313\ : Span4Mux_h
    port map (
            O => \N__33231\,
            I => \N__33180\
        );

    \I__6312\ : Span4Mux_v
    port map (
            O => \N__33224\,
            I => \N__33180\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__33217\,
            I => \N__33177\
        );

    \I__6310\ : Span4Mux_h
    port map (
            O => \N__33212\,
            I => \N__33172\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__33207\,
            I => \N__33172\
        );

    \I__6308\ : InMux
    port map (
            O => \N__33206\,
            I => \N__33163\
        );

    \I__6307\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33163\
        );

    \I__6306\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33163\
        );

    \I__6305\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33163\
        );

    \I__6304\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33160\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__33197\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6302\ : Odrv4
    port map (
            O => \N__33188\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6301\ : Odrv4
    port map (
            O => \N__33185\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6300\ : Odrv4
    port map (
            O => \N__33180\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6299\ : Odrv4
    port map (
            O => \N__33177\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6298\ : Odrv4
    port map (
            O => \N__33172\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__33163\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__33160\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6295\ : InMux
    port map (
            O => \N__33143\,
            I => \N__33133\
        );

    \I__6294\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33124\
        );

    \I__6293\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33119\
        );

    \I__6292\ : InMux
    port map (
            O => \N__33140\,
            I => \N__33114\
        );

    \I__6291\ : InMux
    port map (
            O => \N__33139\,
            I => \N__33114\
        );

    \I__6290\ : InMux
    port map (
            O => \N__33138\,
            I => \N__33107\
        );

    \I__6289\ : InMux
    port map (
            O => \N__33137\,
            I => \N__33107\
        );

    \I__6288\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33107\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__33133\,
            I => \N__33104\
        );

    \I__6286\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33099\
        );

    \I__6285\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33099\
        );

    \I__6284\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33094\
        );

    \I__6283\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33094\
        );

    \I__6282\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33091\
        );

    \I__6281\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33086\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__33124\,
            I => \N__33083\
        );

    \I__6279\ : InMux
    port map (
            O => \N__33123\,
            I => \N__33078\
        );

    \I__6278\ : InMux
    port map (
            O => \N__33122\,
            I => \N__33078\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__33119\,
            I => \N__33072\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__33114\,
            I => \N__33069\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__33107\,
            I => \N__33060\
        );

    \I__6274\ : Span4Mux_h
    port map (
            O => \N__33104\,
            I => \N__33060\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__33099\,
            I => \N__33060\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__33094\,
            I => \N__33060\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__33091\,
            I => \N__33055\
        );

    \I__6270\ : InMux
    port map (
            O => \N__33090\,
            I => \N__33050\
        );

    \I__6269\ : InMux
    port map (
            O => \N__33089\,
            I => \N__33050\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__33086\,
            I => \N__33038\
        );

    \I__6267\ : Span4Mux_h
    port map (
            O => \N__33083\,
            I => \N__33033\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__33078\,
            I => \N__33033\
        );

    \I__6265\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33030\
        );

    \I__6264\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33025\
        );

    \I__6263\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33025\
        );

    \I__6262\ : Span4Mux_h
    port map (
            O => \N__33072\,
            I => \N__33018\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__33069\,
            I => \N__33018\
        );

    \I__6260\ : Span4Mux_v
    port map (
            O => \N__33060\,
            I => \N__33018\
        );

    \I__6259\ : InMux
    port map (
            O => \N__33059\,
            I => \N__33013\
        );

    \I__6258\ : InMux
    port map (
            O => \N__33058\,
            I => \N__33013\
        );

    \I__6257\ : Span4Mux_h
    port map (
            O => \N__33055\,
            I => \N__33008\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__33050\,
            I => \N__33008\
        );

    \I__6255\ : InMux
    port map (
            O => \N__33049\,
            I => \N__32999\
        );

    \I__6254\ : InMux
    port map (
            O => \N__33048\,
            I => \N__32999\
        );

    \I__6253\ : InMux
    port map (
            O => \N__33047\,
            I => \N__32999\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33046\,
            I => \N__32999\
        );

    \I__6251\ : InMux
    port map (
            O => \N__33045\,
            I => \N__32988\
        );

    \I__6250\ : InMux
    port map (
            O => \N__33044\,
            I => \N__32988\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33043\,
            I => \N__32988\
        );

    \I__6248\ : InMux
    port map (
            O => \N__33042\,
            I => \N__32988\
        );

    \I__6247\ : InMux
    port map (
            O => \N__33041\,
            I => \N__32988\
        );

    \I__6246\ : Odrv4
    port map (
            O => \N__33038\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__33033\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__33030\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__33025\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__6242\ : Odrv4
    port map (
            O => \N__33018\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__33013\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__33008\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__32999\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__32988\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__6237\ : InMux
    port map (
            O => \N__32969\,
            I => \N__32964\
        );

    \I__6236\ : InMux
    port map (
            O => \N__32968\,
            I => \N__32961\
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__32967\,
            I => \N__32958\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__32964\,
            I => \N__32955\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__32961\,
            I => \N__32952\
        );

    \I__6232\ : InMux
    port map (
            O => \N__32958\,
            I => \N__32949\
        );

    \I__6231\ : Sp12to4
    port map (
            O => \N__32955\,
            I => \N__32946\
        );

    \I__6230\ : Span4Mux_h
    port map (
            O => \N__32952\,
            I => \N__32943\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__32949\,
            I => measured_delay_hc_22
        );

    \I__6228\ : Odrv12
    port map (
            O => \N__32946\,
            I => measured_delay_hc_22
        );

    \I__6227\ : Odrv4
    port map (
            O => \N__32943\,
            I => measured_delay_hc_22
        );

    \I__6226\ : CascadeMux
    port map (
            O => \N__32936\,
            I => \N__32931\
        );

    \I__6225\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32928\
        );

    \I__6224\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32924\
        );

    \I__6223\ : InMux
    port map (
            O => \N__32931\,
            I => \N__32921\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__32928\,
            I => \N__32917\
        );

    \I__6221\ : InMux
    port map (
            O => \N__32927\,
            I => \N__32914\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__32924\,
            I => \N__32909\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__32921\,
            I => \N__32909\
        );

    \I__6218\ : CascadeMux
    port map (
            O => \N__32920\,
            I => \N__32906\
        );

    \I__6217\ : Span4Mux_v
    port map (
            O => \N__32917\,
            I => \N__32899\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__32914\,
            I => \N__32899\
        );

    \I__6215\ : Span4Mux_h
    port map (
            O => \N__32909\,
            I => \N__32899\
        );

    \I__6214\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32896\
        );

    \I__6213\ : Span4Mux_h
    port map (
            O => \N__32899\,
            I => \N__32893\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__32896\,
            I => measured_delay_hc_16
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__32893\,
            I => measured_delay_hc_16
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__32888\,
            I => \N__32885\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32885\,
            I => \N__32882\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__32882\,
            I => \N__32879\
        );

    \I__6207\ : Odrv4
    port map (
            O => \N__32879\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32876\,
            I => \N__32872\
        );

    \I__6205\ : InMux
    port map (
            O => \N__32875\,
            I => \N__32867\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__32872\,
            I => \N__32863\
        );

    \I__6203\ : InMux
    port map (
            O => \N__32871\,
            I => \N__32858\
        );

    \I__6202\ : InMux
    port map (
            O => \N__32870\,
            I => \N__32858\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__32867\,
            I => \N__32855\
        );

    \I__6200\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32852\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__32863\,
            I => \N__32847\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__32858\,
            I => \N__32847\
        );

    \I__6197\ : Span12Mux_s11_h
    port map (
            O => \N__32855\,
            I => \N__32844\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__32852\,
            I => \N__32841\
        );

    \I__6195\ : Span4Mux_v
    port map (
            O => \N__32847\,
            I => \N__32838\
        );

    \I__6194\ : Odrv12
    port map (
            O => \N__32844\,
            I => measured_delay_hc_1
        );

    \I__6193\ : Odrv4
    port map (
            O => \N__32841\,
            I => measured_delay_hc_1
        );

    \I__6192\ : Odrv4
    port map (
            O => \N__32838\,
            I => measured_delay_hc_1
        );

    \I__6191\ : CascadeMux
    port map (
            O => \N__32831\,
            I => \N__32828\
        );

    \I__6190\ : InMux
    port map (
            O => \N__32828\,
            I => \N__32825\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__32825\,
            I => \N__32822\
        );

    \I__6188\ : Odrv12
    port map (
            O => \N__32822\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__6187\ : InMux
    port map (
            O => \N__32819\,
            I => \N__32811\
        );

    \I__6186\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32811\
        );

    \I__6185\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32806\
        );

    \I__6184\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32806\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__32811\,
            I => \N__32803\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__32806\,
            I => \N__32800\
        );

    \I__6181\ : Odrv4
    port map (
            O => \N__32803\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__6180\ : Odrv12
    port map (
            O => \N__32800\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__6179\ : InMux
    port map (
            O => \N__32795\,
            I => \N__32791\
        );

    \I__6178\ : InMux
    port map (
            O => \N__32794\,
            I => \N__32785\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__32791\,
            I => \N__32782\
        );

    \I__6176\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32779\
        );

    \I__6175\ : CascadeMux
    port map (
            O => \N__32789\,
            I => \N__32776\
        );

    \I__6174\ : CascadeMux
    port map (
            O => \N__32788\,
            I => \N__32773\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__32785\,
            I => \N__32770\
        );

    \I__6172\ : Span4Mux_h
    port map (
            O => \N__32782\,
            I => \N__32767\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__32779\,
            I => \N__32764\
        );

    \I__6170\ : InMux
    port map (
            O => \N__32776\,
            I => \N__32759\
        );

    \I__6169\ : InMux
    port map (
            O => \N__32773\,
            I => \N__32759\
        );

    \I__6168\ : Span4Mux_v
    port map (
            O => \N__32770\,
            I => \N__32756\
        );

    \I__6167\ : Span4Mux_v
    port map (
            O => \N__32767\,
            I => \N__32749\
        );

    \I__6166\ : Span4Mux_h
    port map (
            O => \N__32764\,
            I => \N__32749\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__32759\,
            I => \N__32749\
        );

    \I__6164\ : Odrv4
    port map (
            O => \N__32756\,
            I => measured_delay_hc_3
        );

    \I__6163\ : Odrv4
    port map (
            O => \N__32749\,
            I => measured_delay_hc_3
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__32744\,
            I => \N__32741\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32738\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__32738\,
            I => \N__32735\
        );

    \I__6159\ : Odrv12
    port map (
            O => \N__32735\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__6158\ : InMux
    port map (
            O => \N__32732\,
            I => \N__32729\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__32729\,
            I => \N__32726\
        );

    \I__6156\ : Span4Mux_v
    port map (
            O => \N__32726\,
            I => \N__32720\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32725\,
            I => \N__32717\
        );

    \I__6154\ : InMux
    port map (
            O => \N__32724\,
            I => \N__32713\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32710\
        );

    \I__6152\ : Sp12to4
    port map (
            O => \N__32720\,
            I => \N__32705\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__32717\,
            I => \N__32705\
        );

    \I__6150\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32702\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__32713\,
            I => measured_delay_hc_7
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__32710\,
            I => measured_delay_hc_7
        );

    \I__6147\ : Odrv12
    port map (
            O => \N__32705\,
            I => measured_delay_hc_7
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__32702\,
            I => measured_delay_hc_7
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__32693\,
            I => \N__32690\
        );

    \I__6144\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32687\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__32687\,
            I => \N__32684\
        );

    \I__6142\ : Span4Mux_v
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__6141\ : Odrv4
    port map (
            O => \N__32681\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32675\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__32675\,
            I => \N__32671\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32667\
        );

    \I__6137\ : Span4Mux_h
    port map (
            O => \N__32671\,
            I => \N__32663\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32660\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__32667\,
            I => \N__32656\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32653\
        );

    \I__6133\ : Span4Mux_v
    port map (
            O => \N__32663\,
            I => \N__32650\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32660\,
            I => \N__32647\
        );

    \I__6131\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32644\
        );

    \I__6130\ : Span4Mux_h
    port map (
            O => \N__32656\,
            I => \N__32639\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__32653\,
            I => \N__32639\
        );

    \I__6128\ : Span4Mux_h
    port map (
            O => \N__32650\,
            I => \N__32636\
        );

    \I__6127\ : Span4Mux_v
    port map (
            O => \N__32647\,
            I => \N__32631\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__32644\,
            I => \N__32631\
        );

    \I__6125\ : Span4Mux_h
    port map (
            O => \N__32639\,
            I => \N__32628\
        );

    \I__6124\ : Odrv4
    port map (
            O => \N__32636\,
            I => measured_delay_hc_8
        );

    \I__6123\ : Odrv4
    port map (
            O => \N__32631\,
            I => measured_delay_hc_8
        );

    \I__6122\ : Odrv4
    port map (
            O => \N__32628\,
            I => measured_delay_hc_8
        );

    \I__6121\ : CascadeMux
    port map (
            O => \N__32621\,
            I => \N__32618\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32618\,
            I => \N__32615\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__32615\,
            I => \N__32612\
        );

    \I__6118\ : Odrv12
    port map (
            O => \N__32612\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__6117\ : CascadeMux
    port map (
            O => \N__32609\,
            I => \N__32606\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32603\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__32603\,
            I => \N__32600\
        );

    \I__6114\ : Span4Mux_h
    port map (
            O => \N__32600\,
            I => \N__32597\
        );

    \I__6113\ : Odrv4
    port map (
            O => \N__32597\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__6112\ : CascadeMux
    port map (
            O => \N__32594\,
            I => \N__32591\
        );

    \I__6111\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32588\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__32588\,
            I => \N__32585\
        );

    \I__6109\ : Span4Mux_h
    port map (
            O => \N__32585\,
            I => \N__32582\
        );

    \I__6108\ : Odrv4
    port map (
            O => \N__32582\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__6107\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32576\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__32576\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13\
        );

    \I__6105\ : CascadeMux
    port map (
            O => \N__32573\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\
        );

    \I__6104\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32566\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32562\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__32566\,
            I => \N__32559\
        );

    \I__6101\ : InMux
    port map (
            O => \N__32565\,
            I => \N__32555\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__32562\,
            I => \N__32552\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__32559\,
            I => \N__32549\
        );

    \I__6098\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32546\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__32555\,
            I => measured_delay_hc_0
        );

    \I__6096\ : Odrv12
    port map (
            O => \N__32552\,
            I => measured_delay_hc_0
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__32549\,
            I => measured_delay_hc_0
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__32546\,
            I => measured_delay_hc_0
        );

    \I__6093\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32534\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__32534\,
            I => \N__32531\
        );

    \I__6091\ : Odrv12
    port map (
            O => \N__32531\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_0\
        );

    \I__6090\ : InMux
    port map (
            O => \N__32528\,
            I => \N__32525\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__32525\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32518\
        );

    \I__6087\ : InMux
    port map (
            O => \N__32521\,
            I => \N__32515\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__32518\,
            I => \N__32512\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__32515\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6084\ : Odrv4
    port map (
            O => \N__32512\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6083\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32504\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__32504\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__6081\ : InMux
    port map (
            O => \N__32501\,
            I => \N__32497\
        );

    \I__6080\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32494\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__32497\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__32494\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32489\,
            I => \N__32486\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__32486\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32483\,
            I => \N__32479\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32482\,
            I => \N__32476\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__32479\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32476\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__6071\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32468\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__32468\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__6069\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32461\
        );

    \I__6068\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32458\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__32461\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__32458\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__6065\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32450\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__32450\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__6063\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32443\
        );

    \I__6062\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32440\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__32443\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__32440\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__6059\ : InMux
    port map (
            O => \N__32435\,
            I => \N__32432\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__32432\,
            I => \N__32427\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32431\,
            I => \N__32422\
        );

    \I__6056\ : InMux
    port map (
            O => \N__32430\,
            I => \N__32419\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__32427\,
            I => \N__32416\
        );

    \I__6054\ : InMux
    port map (
            O => \N__32426\,
            I => \N__32413\
        );

    \I__6053\ : InMux
    port map (
            O => \N__32425\,
            I => \N__32410\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__32422\,
            I => \N__32407\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__32419\,
            I => \N__32404\
        );

    \I__6050\ : Span4Mux_v
    port map (
            O => \N__32416\,
            I => \N__32401\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__32413\,
            I => \N__32398\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__32410\,
            I => \N__32395\
        );

    \I__6047\ : Span4Mux_h
    port map (
            O => \N__32407\,
            I => \N__32390\
        );

    \I__6046\ : Span4Mux_h
    port map (
            O => \N__32404\,
            I => \N__32390\
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__32401\,
            I => measured_delay_hc_4
        );

    \I__6044\ : Odrv12
    port map (
            O => \N__32398\,
            I => measured_delay_hc_4
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__32395\,
            I => measured_delay_hc_4
        );

    \I__6042\ : Odrv4
    port map (
            O => \N__32390\,
            I => measured_delay_hc_4
        );

    \I__6041\ : CascadeMux
    port map (
            O => \N__32381\,
            I => \N__32378\
        );

    \I__6040\ : InMux
    port map (
            O => \N__32378\,
            I => \N__32375\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__32375\,
            I => \N__32372\
        );

    \I__6038\ : Odrv12
    port map (
            O => \N__32372\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__6037\ : InMux
    port map (
            O => \N__32369\,
            I => \N__32366\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__32366\,
            I => \N__32361\
        );

    \I__6035\ : InMux
    port map (
            O => \N__32365\,
            I => \N__32358\
        );

    \I__6034\ : InMux
    port map (
            O => \N__32364\,
            I => \N__32353\
        );

    \I__6033\ : Span4Mux_v
    port map (
            O => \N__32361\,
            I => \N__32350\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__32358\,
            I => \N__32347\
        );

    \I__6031\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32344\
        );

    \I__6030\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32341\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__32353\,
            I => \N__32338\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__32350\,
            I => measured_delay_hc_5
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__32347\,
            I => measured_delay_hc_5
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__32344\,
            I => measured_delay_hc_5
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__32341\,
            I => measured_delay_hc_5
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__32338\,
            I => measured_delay_hc_5
        );

    \I__6023\ : CascadeMux
    port map (
            O => \N__32327\,
            I => \N__32324\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32321\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__32321\,
            I => \N__32318\
        );

    \I__6020\ : Span4Mux_h
    port map (
            O => \N__32318\,
            I => \N__32315\
        );

    \I__6019\ : Odrv4
    port map (
            O => \N__32315\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__6018\ : CascadeMux
    port map (
            O => \N__32312\,
            I => \N__32309\
        );

    \I__6017\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32306\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__32306\,
            I => \N__32303\
        );

    \I__6015\ : Span4Mux_h
    port map (
            O => \N__32303\,
            I => \N__32300\
        );

    \I__6014\ : Odrv4
    port map (
            O => \N__32300\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__6013\ : CascadeMux
    port map (
            O => \N__32297\,
            I => \N__32294\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32294\,
            I => \N__32291\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__32291\,
            I => \N__32288\
        );

    \I__6010\ : Span4Mux_h
    port map (
            O => \N__32288\,
            I => \N__32285\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__32285\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__6008\ : InMux
    port map (
            O => \N__32282\,
            I => \N__32279\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__32279\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\
        );

    \I__6006\ : InMux
    port map (
            O => \N__32276\,
            I => \N__32273\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__32273\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\
        );

    \I__6004\ : InMux
    port map (
            O => \N__32270\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__6003\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32264\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__6001\ : Span4Mux_h
    port map (
            O => \N__32261\,
            I => \N__32258\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__32258\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__5999\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32252\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__32252\,
            I => \N__32249\
        );

    \I__5997\ : Span4Mux_v
    port map (
            O => \N__32249\,
            I => \N__32246\
        );

    \I__5996\ : Odrv4
    port map (
            O => \N__32246\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__5995\ : InMux
    port map (
            O => \N__32243\,
            I => \N__32240\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__32240\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__5993\ : InMux
    port map (
            O => \N__32237\,
            I => \N__32233\
        );

    \I__5992\ : InMux
    port map (
            O => \N__32236\,
            I => \N__32230\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__32233\,
            I => \N__32227\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__32230\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5989\ : Odrv4
    port map (
            O => \N__32227\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5988\ : InMux
    port map (
            O => \N__32222\,
            I => \N__32219\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__32219\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__5986\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32212\
        );

    \I__5985\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32209\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__32212\,
            I => \N__32206\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__32209\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__32206\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5981\ : InMux
    port map (
            O => \N__32201\,
            I => \N__32198\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__32198\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32195\,
            I => \N__32191\
        );

    \I__5978\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32188\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__32191\,
            I => \N__32185\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__32188\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__32185\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32177\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__32177\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__5972\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32171\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__32171\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__5970\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32165\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__32165\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__5968\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32159\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__32159\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__5966\ : CascadeMux
    port map (
            O => \N__32156\,
            I => \N__32153\
        );

    \I__5965\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32150\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__32150\,
            I => \N__32147\
        );

    \I__5963\ : Span4Mux_h
    port map (
            O => \N__32147\,
            I => \N__32144\
        );

    \I__5962\ : Odrv4
    port map (
            O => \N__32144\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__5961\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32138\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__32138\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__5959\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32132\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__32132\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__5957\ : InMux
    port map (
            O => \N__32129\,
            I => \N__32126\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__32126\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\
        );

    \I__5955\ : CascadeMux
    port map (
            O => \N__32123\,
            I => \N__32120\
        );

    \I__5954\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32117\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__32117\,
            I => \N__32114\
        );

    \I__5952\ : Odrv4
    port map (
            O => \N__32114\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__5951\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32108\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__32108\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\
        );

    \I__5949\ : InMux
    port map (
            O => \N__32105\,
            I => \N__32102\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__32102\,
            I => \N__32098\
        );

    \I__5947\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32095\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__32098\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__32095\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5944\ : InMux
    port map (
            O => \N__32090\,
            I => \N__32087\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__32087\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__5942\ : CascadeMux
    port map (
            O => \N__32084\,
            I => \N__32081\
        );

    \I__5941\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32077\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32074\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__32077\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__32074\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5937\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32066\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__32066\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__5935\ : InMux
    port map (
            O => \N__32063\,
            I => \N__32059\
        );

    \I__5934\ : InMux
    port map (
            O => \N__32062\,
            I => \N__32056\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__32059\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__32056\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5931\ : InMux
    port map (
            O => \N__32051\,
            I => \N__32048\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__32048\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__5929\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32041\
        );

    \I__5928\ : InMux
    port map (
            O => \N__32044\,
            I => \N__32038\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__32041\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__32038\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5925\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32030\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__32030\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__5923\ : CascadeMux
    port map (
            O => \N__32027\,
            I => \N__32024\
        );

    \I__5922\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32021\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32021\,
            I => \N__32018\
        );

    \I__5920\ : Span4Mux_h
    port map (
            O => \N__32018\,
            I => \N__32015\
        );

    \I__5919\ : Odrv4
    port map (
            O => \N__32015\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ1Z_6\
        );

    \I__5918\ : InMux
    port map (
            O => \N__32012\,
            I => \N__32008\
        );

    \I__5917\ : InMux
    port map (
            O => \N__32011\,
            I => \N__32005\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__32008\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__32005\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5914\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31997\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__31997\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__5912\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31990\
        );

    \I__5911\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31987\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__31990\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__31987\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5908\ : InMux
    port map (
            O => \N__31982\,
            I => \N__31979\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__31979\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__5906\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31973\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__31973\,
            I => \N__31969\
        );

    \I__5904\ : InMux
    port map (
            O => \N__31972\,
            I => \N__31966\
        );

    \I__5903\ : Odrv4
    port map (
            O => \N__31969\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__31966\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5901\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31958\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__31958\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__5899\ : CascadeMux
    port map (
            O => \N__31955\,
            I => \N__31952\
        );

    \I__5898\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31949\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__31949\,
            I => \N__31946\
        );

    \I__5896\ : Span4Mux_h
    port map (
            O => \N__31946\,
            I => \N__31943\
        );

    \I__5895\ : Odrv4
    port map (
            O => \N__31943\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__5894\ : InMux
    port map (
            O => \N__31940\,
            I => \N__31937\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__31937\,
            I => \N__31933\
        );

    \I__5892\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31930\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__31933\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__31930\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5889\ : InMux
    port map (
            O => \N__31925\,
            I => \N__31922\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__31922\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__5887\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31913\
        );

    \I__5886\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31909\
        );

    \I__5885\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31906\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__31916\,
            I => \N__31903\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__31913\,
            I => \N__31900\
        );

    \I__5882\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31897\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__31909\,
            I => \N__31894\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__31906\,
            I => \N__31891\
        );

    \I__5879\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31888\
        );

    \I__5878\ : Span4Mux_v
    port map (
            O => \N__31900\,
            I => \N__31885\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__31897\,
            I => \N__31882\
        );

    \I__5876\ : Span4Mux_v
    port map (
            O => \N__31894\,
            I => \N__31877\
        );

    \I__5875\ : Span4Mux_v
    port map (
            O => \N__31891\,
            I => \N__31877\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__31888\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__31885\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__31882\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__5871\ : Odrv4
    port map (
            O => \N__31877\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__31868\,
            I => \N__31865\
        );

    \I__5869\ : InMux
    port map (
            O => \N__31865\,
            I => \N__31862\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__31862\,
            I => \N__31859\
        );

    \I__5867\ : Odrv4
    port map (
            O => \N__31859\,
            I => \current_shift_inst.PI_CTRL.integrator_i_11\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__31856\,
            I => \N__31851\
        );

    \I__5865\ : CascadeMux
    port map (
            O => \N__31855\,
            I => \N__31848\
        );

    \I__5864\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31843\
        );

    \I__5863\ : InMux
    port map (
            O => \N__31851\,
            I => \N__31840\
        );

    \I__5862\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31837\
        );

    \I__5861\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31834\
        );

    \I__5860\ : InMux
    port map (
            O => \N__31846\,
            I => \N__31831\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__31843\,
            I => \N__31828\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__31840\,
            I => \N__31825\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__31837\,
            I => \N__31822\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__31834\,
            I => \N__31819\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__31831\,
            I => \N__31814\
        );

    \I__5854\ : Span4Mux_h
    port map (
            O => \N__31828\,
            I => \N__31814\
        );

    \I__5853\ : Span4Mux_h
    port map (
            O => \N__31825\,
            I => \N__31809\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__31822\,
            I => \N__31809\
        );

    \I__5851\ : Span4Mux_h
    port map (
            O => \N__31819\,
            I => \N__31806\
        );

    \I__5850\ : Span4Mux_v
    port map (
            O => \N__31814\,
            I => \N__31803\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__31809\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__31806\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5847\ : Odrv4
    port map (
            O => \N__31803\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5846\ : CascadeMux
    port map (
            O => \N__31796\,
            I => \N__31792\
        );

    \I__5845\ : InMux
    port map (
            O => \N__31795\,
            I => \N__31789\
        );

    \I__5844\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31786\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__31789\,
            I => \N__31781\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__31786\,
            I => \N__31778\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__31785\,
            I => \N__31775\
        );

    \I__5840\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31771\
        );

    \I__5839\ : Span4Mux_v
    port map (
            O => \N__31781\,
            I => \N__31768\
        );

    \I__5838\ : Span4Mux_v
    port map (
            O => \N__31778\,
            I => \N__31765\
        );

    \I__5837\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31762\
        );

    \I__5836\ : InMux
    port map (
            O => \N__31774\,
            I => \N__31759\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__31771\,
            I => \N__31756\
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__31768\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__5833\ : Odrv4
    port map (
            O => \N__31765\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__31762\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__31759\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__5830\ : Odrv12
    port map (
            O => \N__31756\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__5829\ : CascadeMux
    port map (
            O => \N__31745\,
            I => \N__31741\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__31744\,
            I => \N__31736\
        );

    \I__5827\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31732\
        );

    \I__5826\ : InMux
    port map (
            O => \N__31740\,
            I => \N__31729\
        );

    \I__5825\ : InMux
    port map (
            O => \N__31739\,
            I => \N__31726\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31736\,
            I => \N__31723\
        );

    \I__5823\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31720\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__31732\,
            I => \N__31717\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__31729\,
            I => \N__31714\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__31726\,
            I => \N__31711\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__31723\,
            I => \N__31708\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__31720\,
            I => \N__31705\
        );

    \I__5817\ : Span4Mux_v
    port map (
            O => \N__31717\,
            I => \N__31702\
        );

    \I__5816\ : Span4Mux_h
    port map (
            O => \N__31714\,
            I => \N__31697\
        );

    \I__5815\ : Span4Mux_h
    port map (
            O => \N__31711\,
            I => \N__31697\
        );

    \I__5814\ : Span4Mux_h
    port map (
            O => \N__31708\,
            I => \N__31692\
        );

    \I__5813\ : Span4Mux_v
    port map (
            O => \N__31705\,
            I => \N__31692\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__31702\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5811\ : Odrv4
    port map (
            O => \N__31697\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__31692\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31679\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__31684\,
            I => \N__31675\
        );

    \I__5807\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31670\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31682\,
            I => \N__31670\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__31679\,
            I => \N__31667\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31664\
        );

    \I__5803\ : InMux
    port map (
            O => \N__31675\,
            I => \N__31661\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__31670\,
            I => \N__31658\
        );

    \I__5801\ : Span4Mux_v
    port map (
            O => \N__31667\,
            I => \N__31655\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__31664\,
            I => \N__31652\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__31661\,
            I => \N__31647\
        );

    \I__5798\ : Span4Mux_v
    port map (
            O => \N__31658\,
            I => \N__31647\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__31655\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5796\ : Odrv4
    port map (
            O => \N__31652\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__31647\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5794\ : InMux
    port map (
            O => \N__31640\,
            I => \N__31637\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31637\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\
        );

    \I__5792\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31631\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__31631\,
            I => \N__31627\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31630\,
            I => \N__31624\
        );

    \I__5789\ : Span4Mux_h
    port map (
            O => \N__31627\,
            I => \N__31621\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__31624\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5787\ : Odrv4
    port map (
            O => \N__31621\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__5786\ : CascadeMux
    port map (
            O => \N__31616\,
            I => \N__31612\
        );

    \I__5785\ : InMux
    port map (
            O => \N__31615\,
            I => \N__31608\
        );

    \I__5784\ : InMux
    port map (
            O => \N__31612\,
            I => \N__31605\
        );

    \I__5783\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31602\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__31608\,
            I => \N__31597\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__31605\,
            I => \N__31592\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31602\,
            I => \N__31592\
        );

    \I__5779\ : InMux
    port map (
            O => \N__31601\,
            I => \N__31587\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31587\
        );

    \I__5777\ : Span12Mux_v
    port map (
            O => \N__31597\,
            I => \N__31584\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__31592\,
            I => \N__31581\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__31587\,
            I => \N__31578\
        );

    \I__5774\ : Odrv12
    port map (
            O => \N__31584\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5773\ : Odrv4
    port map (
            O => \N__31581\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__31578\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__31571\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16_cascade_\
        );

    \I__5770\ : InMux
    port map (
            O => \N__31568\,
            I => \N__31565\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__31565\,
            I => \N__31562\
        );

    \I__5768\ : Span4Mux_h
    port map (
            O => \N__31562\,
            I => \N__31559\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__31559\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\
        );

    \I__5766\ : InMux
    port map (
            O => \N__31556\,
            I => \N__31553\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__31553\,
            I => \N__31550\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__31550\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\
        );

    \I__5763\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31543\
        );

    \I__5762\ : InMux
    port map (
            O => \N__31546\,
            I => \N__31540\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__31543\,
            I => \N__31534\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__31540\,
            I => \N__31534\
        );

    \I__5759\ : InMux
    port map (
            O => \N__31539\,
            I => \N__31531\
        );

    \I__5758\ : Span4Mux_h
    port map (
            O => \N__31534\,
            I => \N__31528\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__31531\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__5756\ : Odrv4
    port map (
            O => \N__31528\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31494\
        );

    \I__5754\ : InMux
    port map (
            O => \N__31522\,
            I => \N__31489\
        );

    \I__5753\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31489\
        );

    \I__5752\ : InMux
    port map (
            O => \N__31520\,
            I => \N__31482\
        );

    \I__5751\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31482\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31518\,
            I => \N__31482\
        );

    \I__5749\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31479\
        );

    \I__5748\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31470\
        );

    \I__5747\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31470\
        );

    \I__5746\ : InMux
    port map (
            O => \N__31514\,
            I => \N__31470\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31513\,
            I => \N__31470\
        );

    \I__5744\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31466\
        );

    \I__5743\ : InMux
    port map (
            O => \N__31511\,
            I => \N__31463\
        );

    \I__5742\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31448\
        );

    \I__5741\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31448\
        );

    \I__5740\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31448\
        );

    \I__5739\ : InMux
    port map (
            O => \N__31507\,
            I => \N__31448\
        );

    \I__5738\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31448\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31448\
        );

    \I__5736\ : InMux
    port map (
            O => \N__31504\,
            I => \N__31448\
        );

    \I__5735\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31433\
        );

    \I__5734\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31433\
        );

    \I__5733\ : InMux
    port map (
            O => \N__31501\,
            I => \N__31433\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31500\,
            I => \N__31433\
        );

    \I__5731\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31433\
        );

    \I__5730\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31433\
        );

    \I__5729\ : InMux
    port map (
            O => \N__31497\,
            I => \N__31433\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__31494\,
            I => \N__31418\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__31489\,
            I => \N__31415\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__31482\,
            I => \N__31408\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__31479\,
            I => \N__31408\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__31470\,
            I => \N__31408\
        );

    \I__5723\ : InMux
    port map (
            O => \N__31469\,
            I => \N__31405\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__31466\,
            I => \N__31402\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__31463\,
            I => \N__31384\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__31448\,
            I => \N__31384\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__31433\,
            I => \N__31384\
        );

    \I__5718\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31375\
        );

    \I__5717\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31375\
        );

    \I__5716\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31375\
        );

    \I__5715\ : InMux
    port map (
            O => \N__31429\,
            I => \N__31375\
        );

    \I__5714\ : InMux
    port map (
            O => \N__31428\,
            I => \N__31372\
        );

    \I__5713\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31357\
        );

    \I__5712\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31357\
        );

    \I__5711\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31357\
        );

    \I__5710\ : InMux
    port map (
            O => \N__31424\,
            I => \N__31357\
        );

    \I__5709\ : InMux
    port map (
            O => \N__31423\,
            I => \N__31357\
        );

    \I__5708\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31357\
        );

    \I__5707\ : InMux
    port map (
            O => \N__31421\,
            I => \N__31357\
        );

    \I__5706\ : Span4Mux_v
    port map (
            O => \N__31418\,
            I => \N__31352\
        );

    \I__5705\ : Span4Mux_v
    port map (
            O => \N__31415\,
            I => \N__31352\
        );

    \I__5704\ : Span4Mux_h
    port map (
            O => \N__31408\,
            I => \N__31349\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__31405\,
            I => \N__31344\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__31402\,
            I => \N__31344\
        );

    \I__5701\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31329\
        );

    \I__5700\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31329\
        );

    \I__5699\ : InMux
    port map (
            O => \N__31399\,
            I => \N__31329\
        );

    \I__5698\ : InMux
    port map (
            O => \N__31398\,
            I => \N__31329\
        );

    \I__5697\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31329\
        );

    \I__5696\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31329\
        );

    \I__5695\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31329\
        );

    \I__5694\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31320\
        );

    \I__5693\ : InMux
    port map (
            O => \N__31393\,
            I => \N__31320\
        );

    \I__5692\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31320\
        );

    \I__5691\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31320\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__31384\,
            I => \N__31315\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__31375\,
            I => \N__31315\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__31372\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__31357\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5686\ : Odrv4
    port map (
            O => \N__31352\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__31349\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__31344\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__31329\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__31320\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5681\ : Odrv4
    port map (
            O => \N__31315\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5680\ : InMux
    port map (
            O => \N__31298\,
            I => \N__31295\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__31295\,
            I => \N__31290\
        );

    \I__5678\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31287\
        );

    \I__5677\ : InMux
    port map (
            O => \N__31293\,
            I => \N__31284\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__31290\,
            I => \N__31281\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__31287\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__31284\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__5673\ : Odrv4
    port map (
            O => \N__31281\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__5672\ : InMux
    port map (
            O => \N__31274\,
            I => \N__31271\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__31271\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__31268\,
            I => \N__31264\
        );

    \I__5669\ : InMux
    port map (
            O => \N__31267\,
            I => \N__31261\
        );

    \I__5668\ : InMux
    port map (
            O => \N__31264\,
            I => \N__31257\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__31261\,
            I => \N__31254\
        );

    \I__5666\ : InMux
    port map (
            O => \N__31260\,
            I => \N__31251\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__31257\,
            I => \N__31246\
        );

    \I__5664\ : Span4Mux_h
    port map (
            O => \N__31254\,
            I => \N__31243\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__31251\,
            I => \N__31240\
        );

    \I__5662\ : InMux
    port map (
            O => \N__31250\,
            I => \N__31235\
        );

    \I__5661\ : InMux
    port map (
            O => \N__31249\,
            I => \N__31235\
        );

    \I__5660\ : Odrv12
    port map (
            O => \N__31246\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5659\ : Odrv4
    port map (
            O => \N__31243\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__31240\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__31235\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5656\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31223\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__31223\,
            I => \N__31220\
        );

    \I__5654\ : Odrv4
    port map (
            O => \N__31220\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\
        );

    \I__5653\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31214\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__31214\,
            I => \N__31211\
        );

    \I__5651\ : Span4Mux_h
    port map (
            O => \N__31211\,
            I => \N__31208\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__31208\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\
        );

    \I__5649\ : InMux
    port map (
            O => \N__31205\,
            I => \N__31201\
        );

    \I__5648\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31198\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__31201\,
            I => \N__31195\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__31198\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5645\ : Odrv4
    port map (
            O => \N__31195\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__5644\ : InMux
    port map (
            O => \N__31190\,
            I => \N__31186\
        );

    \I__5643\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31182\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__31186\,
            I => \N__31178\
        );

    \I__5641\ : InMux
    port map (
            O => \N__31185\,
            I => \N__31174\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__31182\,
            I => \N__31171\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31181\,
            I => \N__31168\
        );

    \I__5638\ : Span4Mux_h
    port map (
            O => \N__31178\,
            I => \N__31165\
        );

    \I__5637\ : InMux
    port map (
            O => \N__31177\,
            I => \N__31162\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__31174\,
            I => \N__31159\
        );

    \I__5635\ : Span12Mux_v
    port map (
            O => \N__31171\,
            I => \N__31154\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__31154\
        );

    \I__5633\ : Odrv4
    port map (
            O => \N__31165\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__31162\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__5631\ : Odrv4
    port map (
            O => \N__31159\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__5630\ : Odrv12
    port map (
            O => \N__31154\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__5629\ : CascadeMux
    port map (
            O => \N__31145\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18_cascade_\
        );

    \I__5628\ : InMux
    port map (
            O => \N__31142\,
            I => \N__31139\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__31139\,
            I => \N__31136\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__31136\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\
        );

    \I__5625\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31130\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__31130\,
            I => \N__31127\
        );

    \I__5623\ : Span4Mux_h
    port map (
            O => \N__31127\,
            I => \N__31124\
        );

    \I__5622\ : Odrv4
    port map (
            O => \N__31124\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\
        );

    \I__5621\ : InMux
    port map (
            O => \N__31121\,
            I => \N__31118\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__31118\,
            I => \N__31113\
        );

    \I__5619\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31110\
        );

    \I__5618\ : InMux
    port map (
            O => \N__31116\,
            I => \N__31107\
        );

    \I__5617\ : Span4Mux_v
    port map (
            O => \N__31113\,
            I => \N__31104\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__31110\,
            I => \N__31101\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__31107\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__31104\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5613\ : Odrv4
    port map (
            O => \N__31101\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__5612\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31090\
        );

    \I__5611\ : InMux
    port map (
            O => \N__31093\,
            I => \N__31087\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__31090\,
            I => \N__31081\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__31087\,
            I => \N__31081\
        );

    \I__5608\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31078\
        );

    \I__5607\ : Span4Mux_v
    port map (
            O => \N__31081\,
            I => \N__31075\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__31078\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__31075\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__5604\ : InMux
    port map (
            O => \N__31070\,
            I => \N__31067\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__31067\,
            I => \N__31064\
        );

    \I__5602\ : Span4Mux_v
    port map (
            O => \N__31064\,
            I => \N__31059\
        );

    \I__5601\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31056\
        );

    \I__5600\ : InMux
    port map (
            O => \N__31062\,
            I => \N__31053\
        );

    \I__5599\ : Span4Mux_v
    port map (
            O => \N__31059\,
            I => \N__31048\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__31056\,
            I => \N__31048\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__31053\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5596\ : Odrv4
    port map (
            O => \N__31048\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__5595\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31039\
        );

    \I__5594\ : InMux
    port map (
            O => \N__31042\,
            I => \N__31036\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__31039\,
            I => \N__31032\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__31036\,
            I => \N__31029\
        );

    \I__5591\ : InMux
    port map (
            O => \N__31035\,
            I => \N__31026\
        );

    \I__5590\ : Span4Mux_h
    port map (
            O => \N__31032\,
            I => \N__31023\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__31029\,
            I => \N__31020\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__31026\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__31023\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__31020\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__5585\ : InMux
    port map (
            O => \N__31013\,
            I => \N__31010\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__31010\,
            I => \N__31007\
        );

    \I__5583\ : Span4Mux_v
    port map (
            O => \N__31007\,
            I => \N__31004\
        );

    \I__5582\ : Odrv4
    port map (
            O => \N__31004\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__31001\,
            I => \N__30998\
        );

    \I__5580\ : InMux
    port map (
            O => \N__30998\,
            I => \N__30995\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__30995\,
            I => \N__30992\
        );

    \I__5578\ : Span4Mux_v
    port map (
            O => \N__30992\,
            I => \N__30989\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__30989\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__5576\ : InMux
    port map (
            O => \N__30986\,
            I => \N__30983\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__30983\,
            I => \N__30980\
        );

    \I__5574\ : Span4Mux_h
    port map (
            O => \N__30980\,
            I => \N__30977\
        );

    \I__5573\ : Span4Mux_h
    port map (
            O => \N__30977\,
            I => \N__30974\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__30974\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__30971\,
            I => \N__30968\
        );

    \I__5570\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30965\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__30965\,
            I => \N__30962\
        );

    \I__5568\ : Span4Mux_h
    port map (
            O => \N__30962\,
            I => \N__30959\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__30959\,
            I => \N__30956\
        );

    \I__5566\ : Odrv4
    port map (
            O => \N__30956\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__5565\ : CascadeMux
    port map (
            O => \N__30953\,
            I => \N__30950\
        );

    \I__5564\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30947\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__30947\,
            I => \N__30944\
        );

    \I__5562\ : Span4Mux_h
    port map (
            O => \N__30944\,
            I => \N__30941\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__30941\,
            I => \current_shift_inst.PI_CTRL.integrator_i_22\
        );

    \I__5560\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30928\
        );

    \I__5559\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30928\
        );

    \I__5558\ : InMux
    port map (
            O => \N__30936\,
            I => \N__30924\
        );

    \I__5557\ : InMux
    port map (
            O => \N__30935\,
            I => \N__30917\
        );

    \I__5556\ : InMux
    port map (
            O => \N__30934\,
            I => \N__30917\
        );

    \I__5555\ : InMux
    port map (
            O => \N__30933\,
            I => \N__30917\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__30928\,
            I => \N__30914\
        );

    \I__5553\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30911\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__30924\,
            I => \delay_measurement_inst.N_299\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__30917\,
            I => \delay_measurement_inst.N_299\
        );

    \I__5550\ : Odrv4
    port map (
            O => \N__30914\,
            I => \delay_measurement_inst.N_299\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__30911\,
            I => \delay_measurement_inst.N_299\
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__30902\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_\
        );

    \I__5547\ : InMux
    port map (
            O => \N__30899\,
            I => \N__30896\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__30896\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5\
        );

    \I__5545\ : CascadeMux
    port map (
            O => \N__30893\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9_cascade_\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__30890\,
            I => \N__30886\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__30889\,
            I => \N__30883\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30886\,
            I => \N__30880\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30877\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__30880\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__30877\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\
        );

    \I__5538\ : CEMux
    port map (
            O => \N__30872\,
            I => \N__30865\
        );

    \I__5537\ : CEMux
    port map (
            O => \N__30871\,
            I => \N__30862\
        );

    \I__5536\ : CEMux
    port map (
            O => \N__30870\,
            I => \N__30859\
        );

    \I__5535\ : CEMux
    port map (
            O => \N__30869\,
            I => \N__30856\
        );

    \I__5534\ : CEMux
    port map (
            O => \N__30868\,
            I => \N__30853\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__30865\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__30862\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__30859\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__30856\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__30853\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__5528\ : CascadeMux
    port map (
            O => \N__30842\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_\
        );

    \I__5527\ : InMux
    port map (
            O => \N__30839\,
            I => \N__30836\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__30836\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\
        );

    \I__5525\ : InMux
    port map (
            O => \N__30833\,
            I => \N__30830\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30830\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5\
        );

    \I__5523\ : InMux
    port map (
            O => \N__30827\,
            I => \N__30824\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__30824\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30818\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__30818\,
            I => \N__30815\
        );

    \I__5519\ : Span4Mux_h
    port map (
            O => \N__30815\,
            I => \N__30812\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__30812\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\
        );

    \I__5517\ : CascadeMux
    port map (
            O => \N__30809\,
            I => \N__30806\
        );

    \I__5516\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30803\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__30803\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\
        );

    \I__5514\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30797\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__30797\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\
        );

    \I__5512\ : CascadeMux
    port map (
            O => \N__30794\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_\
        );

    \I__5511\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30788\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__30788\,
            I => \N__30785\
        );

    \I__5509\ : Odrv4
    port map (
            O => \N__30785\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__30782\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__30779\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6_cascade_\
        );

    \I__5506\ : InMux
    port map (
            O => \N__30776\,
            I => \N__30773\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__30773\,
            I => \delay_measurement_inst.N_42\
        );

    \I__5504\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30767\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__30767\,
            I => \N__30761\
        );

    \I__5502\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30758\
        );

    \I__5501\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30755\
        );

    \I__5500\ : CascadeMux
    port map (
            O => \N__30764\,
            I => \N__30752\
        );

    \I__5499\ : Span4Mux_h
    port map (
            O => \N__30761\,
            I => \N__30749\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__30758\,
            I => \N__30743\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__30755\,
            I => \N__30743\
        );

    \I__5496\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30740\
        );

    \I__5495\ : Span4Mux_h
    port map (
            O => \N__30749\,
            I => \N__30737\
        );

    \I__5494\ : InMux
    port map (
            O => \N__30748\,
            I => \N__30734\
        );

    \I__5493\ : Span4Mux_h
    port map (
            O => \N__30743\,
            I => \N__30731\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__30740\,
            I => \N__30728\
        );

    \I__5491\ : Odrv4
    port map (
            O => \N__30737\,
            I => measured_delay_hc_18
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__30734\,
            I => measured_delay_hc_18
        );

    \I__5489\ : Odrv4
    port map (
            O => \N__30731\,
            I => measured_delay_hc_18
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__30728\,
            I => measured_delay_hc_18
        );

    \I__5487\ : InMux
    port map (
            O => \N__30719\,
            I => \N__30716\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__30716\,
            I => \delay_measurement_inst.N_26\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30713\,
            I => \N__30710\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__30710\,
            I => \N__30707\
        );

    \I__5483\ : Span4Mux_h
    port map (
            O => \N__30707\,
            I => \N__30704\
        );

    \I__5482\ : Span4Mux_v
    port map (
            O => \N__30704\,
            I => \N__30699\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30696\
        );

    \I__5480\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30693\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__30699\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__30696\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__30693\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5476\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30683\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30683\,
            I => \N__30680\
        );

    \I__5474\ : Span4Mux_v
    port map (
            O => \N__30680\,
            I => \N__30674\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30679\,
            I => \N__30669\
        );

    \I__5472\ : InMux
    port map (
            O => \N__30678\,
            I => \N__30669\
        );

    \I__5471\ : InMux
    port map (
            O => \N__30677\,
            I => \N__30666\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__30674\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__30669\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__30666\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5467\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30656\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__30656\,
            I => \N__30653\
        );

    \I__5465\ : Span4Mux_h
    port map (
            O => \N__30653\,
            I => \N__30650\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__30650\,
            I => \delay_measurement_inst.N_27\
        );

    \I__5463\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30644\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__30644\,
            I => \N__30641\
        );

    \I__5461\ : Span4Mux_h
    port map (
            O => \N__30641\,
            I => \N__30637\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30640\,
            I => \N__30634\
        );

    \I__5459\ : Odrv4
    port map (
            O => \N__30637\,
            I => \delay_measurement_inst.elapsed_time_hc_29\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__30634\,
            I => \delay_measurement_inst.elapsed_time_hc_29\
        );

    \I__5457\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30626\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__30626\,
            I => \delay_measurement_inst.N_53\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30619\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30616\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__30619\,
            I => measured_delay_hc_29
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__30616\,
            I => measured_delay_hc_29
        );

    \I__5451\ : InMux
    port map (
            O => \N__30611\,
            I => \N__30608\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__30608\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3\
        );

    \I__5449\ : InMux
    port map (
            O => \N__30605\,
            I => \N__30602\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__30602\,
            I => \delay_measurement_inst.N_54\
        );

    \I__5447\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30595\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30592\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__30595\,
            I => measured_delay_hc_30
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__30592\,
            I => measured_delay_hc_30
        );

    \I__5443\ : InMux
    port map (
            O => \N__30587\,
            I => \N__30584\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__30584\,
            I => \N__30581\
        );

    \I__5441\ : Span4Mux_h
    port map (
            O => \N__30581\,
            I => \N__30578\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__30578\,
            I => delay_hc_input_c
        );

    \I__5439\ : InMux
    port map (
            O => \N__30575\,
            I => \N__30572\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__30572\,
            I => delay_hc_d1
        );

    \I__5437\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30566\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__30566\,
            I => \N__30560\
        );

    \I__5435\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30555\
        );

    \I__5434\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30555\
        );

    \I__5433\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30552\
        );

    \I__5432\ : Span4Mux_h
    port map (
            O => \N__30560\,
            I => \N__30547\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30555\,
            I => \N__30547\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__30552\,
            I => \N__30544\
        );

    \I__5429\ : Span4Mux_v
    port map (
            O => \N__30547\,
            I => \N__30541\
        );

    \I__5428\ : Span4Mux_h
    port map (
            O => \N__30544\,
            I => \N__30538\
        );

    \I__5427\ : Odrv4
    port map (
            O => \N__30541\,
            I => delay_hc_d2
        );

    \I__5426\ : Odrv4
    port map (
            O => \N__30538\,
            I => delay_hc_d2
        );

    \I__5425\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30530\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__30530\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__30527\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30521\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30518\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__30518\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\
        );

    \I__5419\ : InMux
    port map (
            O => \N__30515\,
            I => \N__30512\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__30512\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3\
        );

    \I__5417\ : CascadeMux
    port map (
            O => \N__30509\,
            I => \N__30506\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30506\,
            I => \N__30501\
        );

    \I__5415\ : InMux
    port map (
            O => \N__30505\,
            I => \N__30498\
        );

    \I__5414\ : InMux
    port map (
            O => \N__30504\,
            I => \N__30495\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__30501\,
            I => measured_delay_hc_20
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__30498\,
            I => measured_delay_hc_20
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__30495\,
            I => measured_delay_hc_20
        );

    \I__5410\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30483\
        );

    \I__5409\ : InMux
    port map (
            O => \N__30487\,
            I => \N__30480\
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__30486\,
            I => \N__30477\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__30483\,
            I => \N__30474\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__30480\,
            I => \N__30471\
        );

    \I__5405\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30468\
        );

    \I__5404\ : Span4Mux_h
    port map (
            O => \N__30474\,
            I => \N__30463\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__30471\,
            I => \N__30463\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__30468\,
            I => \N__30460\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__30463\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__5400\ : Odrv4
    port map (
            O => \N__30460\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__30455\,
            I => \delay_measurement_inst.N_29_cascade_\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__30452\,
            I => \N__30448\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__30451\,
            I => \N__30444\
        );

    \I__5396\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30441\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30447\,
            I => \N__30438\
        );

    \I__5394\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30435\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__30441\,
            I => \N__30431\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__30438\,
            I => \N__30426\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__30435\,
            I => \N__30426\
        );

    \I__5390\ : InMux
    port map (
            O => \N__30434\,
            I => \N__30423\
        );

    \I__5389\ : Span4Mux_v
    port map (
            O => \N__30431\,
            I => \N__30419\
        );

    \I__5388\ : Span4Mux_v
    port map (
            O => \N__30426\,
            I => \N__30414\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__30423\,
            I => \N__30414\
        );

    \I__5386\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30411\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__30419\,
            I => \N__30408\
        );

    \I__5384\ : Span4Mux_v
    port map (
            O => \N__30414\,
            I => \N__30405\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__30411\,
            I => measured_delay_hc_6
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__30408\,
            I => measured_delay_hc_6
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__30405\,
            I => measured_delay_hc_6
        );

    \I__5380\ : InMux
    port map (
            O => \N__30398\,
            I => \N__30395\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__30395\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__30392\,
            I => \N__30388\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__30391\,
            I => \N__30384\
        );

    \I__5376\ : InMux
    port map (
            O => \N__30388\,
            I => \N__30381\
        );

    \I__5375\ : CascadeMux
    port map (
            O => \N__30387\,
            I => \N__30378\
        );

    \I__5374\ : InMux
    port map (
            O => \N__30384\,
            I => \N__30375\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__30381\,
            I => \N__30372\
        );

    \I__5372\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30369\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__30375\,
            I => measured_delay_hc_21
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__30372\,
            I => measured_delay_hc_21
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__30369\,
            I => measured_delay_hc_21
        );

    \I__5368\ : InMux
    port map (
            O => \N__30362\,
            I => \N__30358\
        );

    \I__5367\ : CascadeMux
    port map (
            O => \N__30361\,
            I => \N__30354\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__30358\,
            I => \N__30350\
        );

    \I__5365\ : InMux
    port map (
            O => \N__30357\,
            I => \N__30346\
        );

    \I__5364\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30341\
        );

    \I__5363\ : InMux
    port map (
            O => \N__30353\,
            I => \N__30341\
        );

    \I__5362\ : Span4Mux_v
    port map (
            O => \N__30350\,
            I => \N__30338\
        );

    \I__5361\ : InMux
    port map (
            O => \N__30349\,
            I => \N__30335\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__30346\,
            I => \N__30332\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__30341\,
            I => \N__30329\
        );

    \I__5358\ : Span4Mux_h
    port map (
            O => \N__30338\,
            I => \N__30324\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__30335\,
            I => \N__30324\
        );

    \I__5356\ : Span4Mux_h
    port map (
            O => \N__30332\,
            I => \N__30319\
        );

    \I__5355\ : Span4Mux_h
    port map (
            O => \N__30329\,
            I => \N__30319\
        );

    \I__5354\ : Odrv4
    port map (
            O => \N__30324\,
            I => measured_delay_hc_14
        );

    \I__5353\ : Odrv4
    port map (
            O => \N__30319\,
            I => measured_delay_hc_14
        );

    \I__5352\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30311\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__30311\,
            I => \N__30308\
        );

    \I__5350\ : Odrv12
    port map (
            O => \N__30308\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt8\
        );

    \I__5349\ : InMux
    port map (
            O => \N__30305\,
            I => \N__30302\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__30302\,
            I => \N__30299\
        );

    \I__5347\ : Odrv12
    port map (
            O => \N__30299\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__5346\ : CascadeMux
    port map (
            O => \N__30296\,
            I => \N__30292\
        );

    \I__5345\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30289\
        );

    \I__5344\ : InMux
    port map (
            O => \N__30292\,
            I => \N__30286\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__30289\,
            I => \N__30282\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__30286\,
            I => \N__30279\
        );

    \I__5341\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30276\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__30282\,
            I => \N__30273\
        );

    \I__5339\ : Span4Mux_h
    port map (
            O => \N__30279\,
            I => \N__30270\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__30276\,
            I => \N__30267\
        );

    \I__5337\ : Span4Mux_h
    port map (
            O => \N__30273\,
            I => \N__30264\
        );

    \I__5336\ : Span4Mux_v
    port map (
            O => \N__30270\,
            I => \N__30261\
        );

    \I__5335\ : Odrv12
    port map (
            O => \N__30267\,
            I => measured_delay_hc_19
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__30264\,
            I => measured_delay_hc_19
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__30261\,
            I => measured_delay_hc_19
        );

    \I__5332\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30251\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__30251\,
            I => \N__30248\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__30248\,
            I => \N__30245\
        );

    \I__5329\ : Odrv4
    port map (
            O => \N__30245\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__5328\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30239\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__30239\,
            I => \N__30235\
        );

    \I__5326\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30232\
        );

    \I__5325\ : Span4Mux_h
    port map (
            O => \N__30235\,
            I => \N__30224\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__30232\,
            I => \N__30224\
        );

    \I__5323\ : InMux
    port map (
            O => \N__30231\,
            I => \N__30221\
        );

    \I__5322\ : InMux
    port map (
            O => \N__30230\,
            I => \N__30218\
        );

    \I__5321\ : InMux
    port map (
            O => \N__30229\,
            I => \N__30215\
        );

    \I__5320\ : Span4Mux_h
    port map (
            O => \N__30224\,
            I => \N__30212\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__30221\,
            I => \N__30209\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30218\,
            I => measured_delay_hc_17
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__30215\,
            I => measured_delay_hc_17
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__30212\,
            I => measured_delay_hc_17
        );

    \I__5315\ : Odrv12
    port map (
            O => \N__30209\,
            I => measured_delay_hc_17
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__30200\,
            I => \N__30197\
        );

    \I__5313\ : InMux
    port map (
            O => \N__30197\,
            I => \N__30194\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__30194\,
            I => \N__30191\
        );

    \I__5311\ : Odrv12
    port map (
            O => \N__30191\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__5310\ : InMux
    port map (
            O => \N__30188\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__5309\ : InMux
    port map (
            O => \N__30185\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30182\,
            I => \bfn_12_15_0_\
        );

    \I__5307\ : InMux
    port map (
            O => \N__30179\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__5306\ : InMux
    port map (
            O => \N__30176\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__5305\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30170\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__30170\,
            I => \N__30167\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__30164\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__5301\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30158\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__30158\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__5299\ : InMux
    port map (
            O => \N__30155\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__5298\ : CascadeMux
    port map (
            O => \N__30152\,
            I => \N__30149\
        );

    \I__5297\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30146\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__30146\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__5295\ : InMux
    port map (
            O => \N__30143\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__5294\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30137\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__30137\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__5292\ : InMux
    port map (
            O => \N__30134\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__5291\ : CascadeMux
    port map (
            O => \N__30131\,
            I => \N__30128\
        );

    \I__5290\ : InMux
    port map (
            O => \N__30128\,
            I => \N__30125\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__30125\,
            I => \N__30122\
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__30122\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__5287\ : InMux
    port map (
            O => \N__30119\,
            I => \bfn_12_14_0_\
        );

    \I__5286\ : InMux
    port map (
            O => \N__30116\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__5285\ : InMux
    port map (
            O => \N__30113\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__5284\ : InMux
    port map (
            O => \N__30110\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30107\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30104\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__5281\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30098\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__30098\,
            I => \N__30095\
        );

    \I__5279\ : Odrv4
    port map (
            O => \N__30095\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__5278\ : InMux
    port map (
            O => \N__30092\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__30089\,
            I => \N__30086\
        );

    \I__5276\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30083\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__30083\,
            I => \N__30080\
        );

    \I__5274\ : Odrv4
    port map (
            O => \N__30080\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__5273\ : InMux
    port map (
            O => \N__30077\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__5272\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30071\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__30071\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30068\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__5269\ : CascadeMux
    port map (
            O => \N__30065\,
            I => \N__30062\
        );

    \I__5268\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30059\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__30059\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__5266\ : InMux
    port map (
            O => \N__30056\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__5265\ : InMux
    port map (
            O => \N__30053\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__5264\ : InMux
    port map (
            O => \N__30050\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__5263\ : InMux
    port map (
            O => \N__30047\,
            I => \N__30044\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__30044\,
            I => \N__30039\
        );

    \I__5261\ : InMux
    port map (
            O => \N__30043\,
            I => \N__30036\
        );

    \I__5260\ : InMux
    port map (
            O => \N__30042\,
            I => \N__30033\
        );

    \I__5259\ : Span4Mux_v
    port map (
            O => \N__30039\,
            I => \N__30028\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__30036\,
            I => \N__30028\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__30033\,
            I => \N__30025\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__30028\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__30025\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__5254\ : InMux
    port map (
            O => \N__30020\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__5253\ : InMux
    port map (
            O => \N__30017\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__5252\ : InMux
    port map (
            O => \N__30014\,
            I => \N__30010\
        );

    \I__5251\ : InMux
    port map (
            O => \N__30013\,
            I => \N__30007\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__30010\,
            I => \N__30001\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__30007\,
            I => \N__30001\
        );

    \I__5248\ : InMux
    port map (
            O => \N__30006\,
            I => \N__29998\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__30001\,
            I => \N__29995\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__29998\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__5245\ : Odrv4
    port map (
            O => \N__29995\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__29990\,
            I => \N__29987\
        );

    \I__5243\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29984\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__29984\,
            I => \N__29981\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__29981\,
            I => \N__29978\
        );

    \I__5240\ : Span4Mux_h
    port map (
            O => \N__29978\,
            I => \N__29975\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__29975\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__5238\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29967\
        );

    \I__5237\ : InMux
    port map (
            O => \N__29971\,
            I => \N__29964\
        );

    \I__5236\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29961\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__29967\,
            I => \N__29958\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__29964\,
            I => \N__29955\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__29961\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__5232\ : Odrv4
    port map (
            O => \N__29958\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__29955\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__29948\,
            I => \N__29945\
        );

    \I__5229\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29942\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__5227\ : Span4Mux_h
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__5226\ : Odrv4
    port map (
            O => \N__29936\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__5225\ : InMux
    port map (
            O => \N__29933\,
            I => \N__29929\
        );

    \I__5224\ : InMux
    port map (
            O => \N__29932\,
            I => \N__29926\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__29929\,
            I => \N__29923\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__29926\,
            I => \N__29920\
        );

    \I__5221\ : Odrv12
    port map (
            O => \N__29923\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__5220\ : Odrv4
    port map (
            O => \N__29920\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__5219\ : InMux
    port map (
            O => \N__29915\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__5218\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29909\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__29909\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__5216\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29902\
        );

    \I__5215\ : InMux
    port map (
            O => \N__29905\,
            I => \N__29899\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__29902\,
            I => \N__29896\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__29899\,
            I => \N__29893\
        );

    \I__5212\ : Odrv4
    port map (
            O => \N__29896\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__5211\ : Odrv4
    port map (
            O => \N__29893\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__5210\ : InMux
    port map (
            O => \N__29888\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__5209\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29882\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__29882\,
            I => \N__29878\
        );

    \I__5207\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29875\
        );

    \I__5206\ : Span4Mux_v
    port map (
            O => \N__29878\,
            I => \N__29872\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__29875\,
            I => \N__29869\
        );

    \I__5204\ : Odrv4
    port map (
            O => \N__29872\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__29869\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5202\ : InMux
    port map (
            O => \N__29864\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__5201\ : InMux
    port map (
            O => \N__29861\,
            I => \N__29857\
        );

    \I__5200\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29854\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__29857\,
            I => \N__29851\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__29854\,
            I => \N__29847\
        );

    \I__5197\ : Span4Mux_h
    port map (
            O => \N__29851\,
            I => \N__29844\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29850\,
            I => \N__29841\
        );

    \I__5195\ : Odrv12
    port map (
            O => \N__29847\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__29844\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__29841\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5192\ : InMux
    port map (
            O => \N__29834\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__5191\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29828\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29825\
        );

    \I__5189\ : Span4Mux_h
    port map (
            O => \N__29825\,
            I => \N__29822\
        );

    \I__5188\ : Odrv4
    port map (
            O => \N__29822\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__5187\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29815\
        );

    \I__5186\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29811\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__29815\,
            I => \N__29808\
        );

    \I__5184\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29805\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__29811\,
            I => \N__29802\
        );

    \I__5182\ : Span4Mux_h
    port map (
            O => \N__29808\,
            I => \N__29799\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__29805\,
            I => \N__29796\
        );

    \I__5180\ : Odrv12
    port map (
            O => \N__29802\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__29799\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__29796\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__5177\ : InMux
    port map (
            O => \N__29789\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29783\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__29783\,
            I => \N__29780\
        );

    \I__5174\ : Span4Mux_h
    port map (
            O => \N__29780\,
            I => \N__29777\
        );

    \I__5173\ : Span4Mux_h
    port map (
            O => \N__29777\,
            I => \N__29774\
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__29774\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29767\
        );

    \I__5170\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29764\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__29767\,
            I => \N__29761\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__29764\,
            I => \N__29757\
        );

    \I__5167\ : Span4Mux_h
    port map (
            O => \N__29761\,
            I => \N__29754\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29751\
        );

    \I__5165\ : Odrv12
    port map (
            O => \N__29757\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__29754\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__29751\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29744\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__5161\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29737\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29734\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__29737\,
            I => \N__29730\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__29734\,
            I => \N__29727\
        );

    \I__5157\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29724\
        );

    \I__5156\ : Span4Mux_h
    port map (
            O => \N__29730\,
            I => \N__29721\
        );

    \I__5155\ : Span4Mux_h
    port map (
            O => \N__29727\,
            I => \N__29716\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__29724\,
            I => \N__29716\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__29721\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__29716\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29711\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29705\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29702\
        );

    \I__5148\ : Span4Mux_h
    port map (
            O => \N__29702\,
            I => \N__29699\
        );

    \I__5147\ : Odrv4
    port map (
            O => \N__29699\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29696\,
            I => \N__29693\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__29693\,
            I => \N__29688\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29685\
        );

    \I__5143\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29682\
        );

    \I__5142\ : Span4Mux_v
    port map (
            O => \N__29688\,
            I => \N__29675\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29685\,
            I => \N__29675\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__29682\,
            I => \N__29675\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__29675\,
            I => \N__29672\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__29672\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29669\,
            I => \bfn_12_11_0_\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__29666\,
            I => \N__29663\
        );

    \I__5135\ : InMux
    port map (
            O => \N__29663\,
            I => \N__29660\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__29660\,
            I => \N__29657\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__29657\,
            I => \N__29654\
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__29654\,
            I => \current_shift_inst.PI_CTRL.integrator_i_14\
        );

    \I__5131\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29647\
        );

    \I__5130\ : InMux
    port map (
            O => \N__29650\,
            I => \N__29643\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__29647\,
            I => \N__29640\
        );

    \I__5128\ : InMux
    port map (
            O => \N__29646\,
            I => \N__29637\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__29643\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__29640\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29637\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__5124\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29626\
        );

    \I__5123\ : InMux
    port map (
            O => \N__29629\,
            I => \N__29622\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__29626\,
            I => \N__29619\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29616\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__29622\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__29619\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__29616\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__5117\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29605\
        );

    \I__5116\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29601\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__29605\,
            I => \N__29598\
        );

    \I__5114\ : InMux
    port map (
            O => \N__29604\,
            I => \N__29595\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__29601\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__5112\ : Odrv4
    port map (
            O => \N__29598\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__29595\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__5110\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__29585\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__29579\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\
        );

    \I__5106\ : InMux
    port map (
            O => \N__29576\,
            I => \N__29573\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__29573\,
            I => \N__29570\
        );

    \I__5104\ : Span4Mux_v
    port map (
            O => \N__29570\,
            I => \N__29565\
        );

    \I__5103\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29562\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29559\
        );

    \I__5101\ : Span4Mux_v
    port map (
            O => \N__29565\,
            I => \N__29556\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__29562\,
            I => \N__29553\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__29559\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__29556\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__5097\ : Odrv12
    port map (
            O => \N__29553\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__5096\ : InMux
    port map (
            O => \N__29546\,
            I => \N__29543\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__29543\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\
        );

    \I__5094\ : InMux
    port map (
            O => \N__29540\,
            I => \N__29537\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__29537\,
            I => \N__29534\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__29534\,
            I => \N__29531\
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__29531\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\
        );

    \I__5090\ : InMux
    port map (
            O => \N__29528\,
            I => \N__29525\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__29525\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__5088\ : CascadeMux
    port map (
            O => \N__29522\,
            I => \N__29519\
        );

    \I__5087\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29513\
        );

    \I__5086\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29510\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__29517\,
            I => \N__29507\
        );

    \I__5084\ : InMux
    port map (
            O => \N__29516\,
            I => \N__29504\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__29513\,
            I => \N__29498\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__29510\,
            I => \N__29498\
        );

    \I__5081\ : InMux
    port map (
            O => \N__29507\,
            I => \N__29495\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__29504\,
            I => \N__29492\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__29503\,
            I => \N__29489\
        );

    \I__5078\ : Span4Mux_h
    port map (
            O => \N__29498\,
            I => \N__29486\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29483\
        );

    \I__5076\ : Span4Mux_h
    port map (
            O => \N__29492\,
            I => \N__29480\
        );

    \I__5075\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29477\
        );

    \I__5074\ : Span4Mux_v
    port map (
            O => \N__29486\,
            I => \N__29474\
        );

    \I__5073\ : Odrv4
    port map (
            O => \N__29483\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__29480\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__29477\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__29474\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__5069\ : CascadeMux
    port map (
            O => \N__29465\,
            I => \N__29462\
        );

    \I__5068\ : InMux
    port map (
            O => \N__29462\,
            I => \N__29459\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__29459\,
            I => \N__29456\
        );

    \I__5066\ : Span4Mux_v
    port map (
            O => \N__29456\,
            I => \N__29453\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__29453\,
            I => \N__29450\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__29450\,
            I => \current_shift_inst.PI_CTRL.integrator_i_20\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__29447\,
            I => \N__29444\
        );

    \I__5062\ : InMux
    port map (
            O => \N__29444\,
            I => \N__29441\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__29441\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\
        );

    \I__5060\ : InMux
    port map (
            O => \N__29438\,
            I => \N__29435\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__29435\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\
        );

    \I__5058\ : InMux
    port map (
            O => \N__29432\,
            I => \N__29429\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__29429\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\
        );

    \I__5056\ : InMux
    port map (
            O => \N__29426\,
            I => \N__29423\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__29423\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\
        );

    \I__5054\ : InMux
    port map (
            O => \N__29420\,
            I => \N__29417\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__29417\,
            I => \delay_measurement_inst.N_59\
        );

    \I__5052\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29406\
        );

    \I__5051\ : InMux
    port map (
            O => \N__29413\,
            I => \N__29395\
        );

    \I__5050\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29395\
        );

    \I__5049\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29395\
        );

    \I__5048\ : InMux
    port map (
            O => \N__29410\,
            I => \N__29395\
        );

    \I__5047\ : InMux
    port map (
            O => \N__29409\,
            I => \N__29395\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__29406\,
            I => \delay_measurement_inst.N_270\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__29395\,
            I => \delay_measurement_inst.N_270\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__29390\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__29387\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7_cascade_\
        );

    \I__5042\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29381\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__29381\,
            I => \N__29378\
        );

    \I__5040\ : Span4Mux_h
    port map (
            O => \N__29378\,
            I => \N__29375\
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__29375\,
            I => delay_tr_input_c
        );

    \I__5038\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29369\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__29369\,
            I => delay_tr_d1
        );

    \I__5036\ : InMux
    port map (
            O => \N__29366\,
            I => \N__29360\
        );

    \I__5035\ : InMux
    port map (
            O => \N__29365\,
            I => \N__29355\
        );

    \I__5034\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29355\
        );

    \I__5033\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29352\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__29360\,
            I => delay_tr_d2
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__29355\,
            I => delay_tr_d2
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__29352\,
            I => delay_tr_d2
        );

    \I__5029\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29340\
        );

    \I__5028\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29337\
        );

    \I__5027\ : InMux
    port map (
            O => \N__29343\,
            I => \N__29334\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__29340\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__29337\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__29334\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__5023\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29322\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29319\
        );

    \I__5021\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29316\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__29322\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__29319\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__29316\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__5017\ : InMux
    port map (
            O => \N__29309\,
            I => \N__29306\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__29306\,
            I => \N__29302\
        );

    \I__5015\ : InMux
    port map (
            O => \N__29305\,
            I => \N__29299\
        );

    \I__5014\ : Span4Mux_v
    port map (
            O => \N__29302\,
            I => \N__29294\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__29299\,
            I => \N__29294\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__29294\,
            I => \N__29291\
        );

    \I__5011\ : Span4Mux_v
    port map (
            O => \N__29291\,
            I => \N__29288\
        );

    \I__5010\ : Span4Mux_v
    port map (
            O => \N__29288\,
            I => \N__29285\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__29285\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5008\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29279\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29275\
        );

    \I__5006\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29272\
        );

    \I__5005\ : Span4Mux_v
    port map (
            O => \N__29275\,
            I => \N__29268\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__29272\,
            I => \N__29265\
        );

    \I__5003\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29262\
        );

    \I__5002\ : Span4Mux_v
    port map (
            O => \N__29268\,
            I => \N__29259\
        );

    \I__5001\ : Span4Mux_h
    port map (
            O => \N__29265\,
            I => \N__29256\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__29262\,
            I => \N__29253\
        );

    \I__4999\ : Sp12to4
    port map (
            O => \N__29259\,
            I => \N__29250\
        );

    \I__4998\ : Sp12to4
    port map (
            O => \N__29256\,
            I => \N__29245\
        );

    \I__4997\ : Sp12to4
    port map (
            O => \N__29253\,
            I => \N__29245\
        );

    \I__4996\ : Span12Mux_h
    port map (
            O => \N__29250\,
            I => \N__29240\
        );

    \I__4995\ : Span12Mux_v
    port map (
            O => \N__29245\,
            I => \N__29240\
        );

    \I__4994\ : Odrv12
    port map (
            O => \N__29240\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29231\
        );

    \I__4992\ : InMux
    port map (
            O => \N__29236\,
            I => \N__29231\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__29231\,
            I => \N__29228\
        );

    \I__4990\ : Span4Mux_v
    port map (
            O => \N__29228\,
            I => \N__29223\
        );

    \I__4989\ : InMux
    port map (
            O => \N__29227\,
            I => \N__29220\
        );

    \I__4988\ : InMux
    port map (
            O => \N__29226\,
            I => \N__29217\
        );

    \I__4987\ : Span4Mux_h
    port map (
            O => \N__29223\,
            I => \N__29214\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__29220\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__29217\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__29214\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4983\ : CascadeMux
    port map (
            O => \N__29207\,
            I => \N__29204\
        );

    \I__4982\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29200\
        );

    \I__4981\ : InMux
    port map (
            O => \N__29203\,
            I => \N__29197\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__29200\,
            I => \N__29192\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__29197\,
            I => \N__29192\
        );

    \I__4978\ : Odrv12
    port map (
            O => \N__29192\,
            I => measured_delay_hc_25
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__29189\,
            I => \N__29186\
        );

    \I__4976\ : InMux
    port map (
            O => \N__29186\,
            I => \N__29182\
        );

    \I__4975\ : InMux
    port map (
            O => \N__29185\,
            I => \N__29179\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__29182\,
            I => measured_delay_hc_24
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__29179\,
            I => measured_delay_hc_24
        );

    \I__4972\ : CascadeMux
    port map (
            O => \N__29174\,
            I => \N__29171\
        );

    \I__4971\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29167\
        );

    \I__4970\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29164\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__29167\,
            I => \N__29161\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__29164\,
            I => measured_delay_hc_26
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__29161\,
            I => measured_delay_hc_26
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__4965\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29149\
        );

    \I__4964\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29146\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__29149\,
            I => measured_delay_hc_23
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__29146\,
            I => measured_delay_hc_23
        );

    \I__4961\ : InMux
    port map (
            O => \N__29141\,
            I => \N__29138\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__29138\,
            I => \N__29134\
        );

    \I__4959\ : InMux
    port map (
            O => \N__29137\,
            I => \N__29131\
        );

    \I__4958\ : Span4Mux_h
    port map (
            O => \N__29134\,
            I => \N__29128\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__29131\,
            I => measured_delay_hc_28
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__29128\,
            I => measured_delay_hc_28
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__29123\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4_cascade_\
        );

    \I__4954\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29116\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__29119\,
            I => \N__29113\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__29116\,
            I => \N__29110\
        );

    \I__4951\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29107\
        );

    \I__4950\ : Odrv4
    port map (
            O => \N__29110\,
            I => \delay_measurement_inst.elapsed_time_hc_30\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29107\,
            I => \delay_measurement_inst.elapsed_time_hc_30\
        );

    \I__4948\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29099\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__29099\,
            I => \delay_measurement_inst.N_51\
        );

    \I__4946\ : InMux
    port map (
            O => \N__29096\,
            I => \N__29093\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__29093\,
            I => \N__29089\
        );

    \I__4944\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29086\
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__29089\,
            I => measured_delay_hc_27
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__29086\,
            I => measured_delay_hc_27
        );

    \I__4941\ : InMux
    port map (
            O => \N__29081\,
            I => \N__29078\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__29078\,
            I => \delay_measurement_inst.N_25\
        );

    \I__4939\ : IoInMux
    port map (
            O => \N__29075\,
            I => \N__29072\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__29072\,
            I => \delay_measurement_inst.delay_tr_timer.N_304_i\
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__29069\,
            I => \delay_measurement_inst.N_33_cascade_\
        );

    \I__4936\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29063\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__29063\,
            I => \N__29060\
        );

    \I__4934\ : Odrv12
    port map (
            O => \N__29060\,
            I => \delay_measurement_inst.N_38\
        );

    \I__4933\ : InMux
    port map (
            O => \N__29057\,
            I => \N__29054\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__29054\,
            I => \N__29049\
        );

    \I__4931\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29044\
        );

    \I__4930\ : InMux
    port map (
            O => \N__29052\,
            I => \N__29044\
        );

    \I__4929\ : Odrv12
    port map (
            O => \N__29049\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__29044\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__4927\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29036\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__29036\,
            I => \N__29032\
        );

    \I__4925\ : InMux
    port map (
            O => \N__29035\,
            I => \N__29029\
        );

    \I__4924\ : Span4Mux_v
    port map (
            O => \N__29032\,
            I => \N__29026\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__29029\,
            I => \N__29023\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__29026\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__29023\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__4920\ : InMux
    port map (
            O => \N__29018\,
            I => \N__29014\
        );

    \I__4919\ : InMux
    port map (
            O => \N__29017\,
            I => \N__29011\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__29014\,
            I => \N__29008\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__29011\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__29008\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\
        );

    \I__4915\ : CascadeMux
    port map (
            O => \N__29003\,
            I => \N__29000\
        );

    \I__4914\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28997\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__28997\,
            I => \N__28994\
        );

    \I__4912\ : Odrv4
    port map (
            O => \N__28994\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_0\
        );

    \I__4911\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28988\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28985\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__28985\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\
        );

    \I__4908\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28978\
        );

    \I__4907\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28974\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__28978\,
            I => \N__28971\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__28977\,
            I => \N__28968\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__28974\,
            I => \N__28965\
        );

    \I__4903\ : Span4Mux_h
    port map (
            O => \N__28971\,
            I => \N__28962\
        );

    \I__4902\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28959\
        );

    \I__4901\ : Span4Mux_h
    port map (
            O => \N__28965\,
            I => \N__28956\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__28962\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__28959\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__4898\ : Odrv4
    port map (
            O => \N__28956\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__4897\ : CEMux
    port map (
            O => \N__28949\,
            I => \N__28945\
        );

    \I__4896\ : CEMux
    port map (
            O => \N__28948\,
            I => \N__28941\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__28945\,
            I => \N__28937\
        );

    \I__4894\ : CEMux
    port map (
            O => \N__28944\,
            I => \N__28934\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__28941\,
            I => \N__28931\
        );

    \I__4892\ : CEMux
    port map (
            O => \N__28940\,
            I => \N__28928\
        );

    \I__4891\ : Span4Mux_v
    port map (
            O => \N__28937\,
            I => \N__28923\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__28934\,
            I => \N__28923\
        );

    \I__4889\ : Span4Mux_v
    port map (
            O => \N__28931\,
            I => \N__28918\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__28928\,
            I => \N__28918\
        );

    \I__4887\ : Sp12to4
    port map (
            O => \N__28923\,
            I => \N__28915\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__28918\,
            I => \delay_measurement_inst.delay_hc_timer.N_303_i\
        );

    \I__4885\ : Odrv12
    port map (
            O => \N__28915\,
            I => \delay_measurement_inst.delay_hc_timer.N_303_i\
        );

    \I__4884\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28907\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__28907\,
            I => \N__28904\
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__28904\,
            I => \delay_measurement_inst.N_28\
        );

    \I__4881\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28896\
        );

    \I__4880\ : InMux
    port map (
            O => \N__28900\,
            I => \N__28893\
        );

    \I__4879\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28890\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__28896\,
            I => \N__28885\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__28893\,
            I => \N__28885\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__28890\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__4875\ : Odrv12
    port map (
            O => \N__28885\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__4874\ : InMux
    port map (
            O => \N__28880\,
            I => \N__28877\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__28877\,
            I => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\
        );

    \I__4872\ : CascadeMux
    port map (
            O => \N__28874\,
            I => \N__28871\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28871\,
            I => \N__28868\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__28868\,
            I => \N__28865\
        );

    \I__4869\ : Span4Mux_h
    port map (
            O => \N__28865\,
            I => \N__28862\
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__28862\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__28859\,
            I => \N__28856\
        );

    \I__4866\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28853\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__28853\,
            I => \N__28850\
        );

    \I__4864\ : Odrv12
    port map (
            O => \N__28850\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__4863\ : CEMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__28844\,
            I => \N__28839\
        );

    \I__4861\ : CEMux
    port map (
            O => \N__28843\,
            I => \N__28836\
        );

    \I__4860\ : CEMux
    port map (
            O => \N__28842\,
            I => \N__28833\
        );

    \I__4859\ : Span4Mux_h
    port map (
            O => \N__28839\,
            I => \N__28828\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__28836\,
            I => \N__28825\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__28833\,
            I => \N__28822\
        );

    \I__4856\ : CEMux
    port map (
            O => \N__28832\,
            I => \N__28819\
        );

    \I__4855\ : CEMux
    port map (
            O => \N__28831\,
            I => \N__28816\
        );

    \I__4854\ : Span4Mux_v
    port map (
            O => \N__28828\,
            I => \N__28813\
        );

    \I__4853\ : Span4Mux_h
    port map (
            O => \N__28825\,
            I => \N__28810\
        );

    \I__4852\ : Span4Mux_v
    port map (
            O => \N__28822\,
            I => \N__28807\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__28819\,
            I => \N__28802\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__28816\,
            I => \N__28802\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__28813\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__28810\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__28807\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__4846\ : Odrv12
    port map (
            O => \N__28802\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__4845\ : InMux
    port map (
            O => \N__28793\,
            I => \N__28790\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__28790\,
            I => \N__28786\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__28789\,
            I => \N__28783\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__28786\,
            I => \N__28780\
        );

    \I__4841\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28777\
        );

    \I__4840\ : Span4Mux_v
    port map (
            O => \N__28780\,
            I => \N__28774\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__28777\,
            I => \N__28771\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__28774\,
            I => \N__28768\
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__28771\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__28768\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__4835\ : InMux
    port map (
            O => \N__28763\,
            I => \N__28760\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__28760\,
            I => \N__28754\
        );

    \I__4833\ : InMux
    port map (
            O => \N__28759\,
            I => \N__28747\
        );

    \I__4832\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28747\
        );

    \I__4831\ : InMux
    port map (
            O => \N__28757\,
            I => \N__28747\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__28754\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__28747\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__4828\ : InMux
    port map (
            O => \N__28742\,
            I => \N__28739\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__28739\,
            I => \N__28736\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__28736\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\
        );

    \I__4825\ : CascadeMux
    port map (
            O => \N__28733\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28730\,
            I => \N__28726\
        );

    \I__4823\ : InMux
    port map (
            O => \N__28729\,
            I => \N__28722\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__28726\,
            I => \N__28719\
        );

    \I__4821\ : InMux
    port map (
            O => \N__28725\,
            I => \N__28716\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__28722\,
            I => \N__28713\
        );

    \I__4819\ : Span4Mux_v
    port map (
            O => \N__28719\,
            I => \N__28708\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__28716\,
            I => \N__28705\
        );

    \I__4817\ : Span4Mux_h
    port map (
            O => \N__28713\,
            I => \N__28702\
        );

    \I__4816\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28697\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28697\
        );

    \I__4814\ : Odrv4
    port map (
            O => \N__28708\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__28705\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__28702\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__28697\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4810\ : InMux
    port map (
            O => \N__28688\,
            I => \N__28685\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__28685\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\
        );

    \I__4808\ : CascadeMux
    port map (
            O => \N__28682\,
            I => \N__28678\
        );

    \I__4807\ : CascadeMux
    port map (
            O => \N__28681\,
            I => \N__28674\
        );

    \I__4806\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28667\
        );

    \I__4805\ : InMux
    port map (
            O => \N__28677\,
            I => \N__28667\
        );

    \I__4804\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28667\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__28667\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_0_16\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__28664\,
            I => \N__28655\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__28663\,
            I => \N__28651\
        );

    \I__4800\ : CascadeMux
    port map (
            O => \N__28662\,
            I => \N__28647\
        );

    \I__4799\ : CascadeMux
    port map (
            O => \N__28661\,
            I => \N__28643\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__28660\,
            I => \N__28639\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__28659\,
            I => \N__28635\
        );

    \I__4796\ : InMux
    port map (
            O => \N__28658\,
            I => \N__28624\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28624\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28624\
        );

    \I__4793\ : InMux
    port map (
            O => \N__28651\,
            I => \N__28624\
        );

    \I__4792\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28607\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28647\,
            I => \N__28607\
        );

    \I__4790\ : InMux
    port map (
            O => \N__28646\,
            I => \N__28607\
        );

    \I__4789\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28607\
        );

    \I__4788\ : InMux
    port map (
            O => \N__28642\,
            I => \N__28607\
        );

    \I__4787\ : InMux
    port map (
            O => \N__28639\,
            I => \N__28607\
        );

    \I__4786\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28607\
        );

    \I__4785\ : InMux
    port map (
            O => \N__28635\,
            I => \N__28607\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__28634\,
            I => \N__28603\
        );

    \I__4783\ : CascadeMux
    port map (
            O => \N__28633\,
            I => \N__28599\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__28624\,
            I => \N__28594\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__28607\,
            I => \N__28594\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28585\
        );

    \I__4779\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28585\
        );

    \I__4778\ : InMux
    port map (
            O => \N__28602\,
            I => \N__28585\
        );

    \I__4777\ : InMux
    port map (
            O => \N__28599\,
            I => \N__28585\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__28594\,
            I => \N__28580\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__28585\,
            I => \N__28580\
        );

    \I__4774\ : Span4Mux_h
    port map (
            O => \N__28580\,
            I => \N__28577\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__28577\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__4772\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28570\
        );

    \I__4771\ : InMux
    port map (
            O => \N__28573\,
            I => \N__28566\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__28570\,
            I => \N__28563\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28569\,
            I => \N__28560\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__28566\,
            I => \N__28557\
        );

    \I__4767\ : Span4Mux_v
    port map (
            O => \N__28563\,
            I => \N__28554\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28560\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__28557\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__28554\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28542\
        );

    \I__4762\ : InMux
    port map (
            O => \N__28546\,
            I => \N__28539\
        );

    \I__4761\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28536\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__28542\,
            I => \N__28533\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28530\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__28536\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__28533\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__4756\ : Odrv12
    port map (
            O => \N__28530\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__4755\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28519\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28516\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__28519\,
            I => \N__28510\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28516\,
            I => \N__28510\
        );

    \I__4751\ : InMux
    port map (
            O => \N__28515\,
            I => \N__28507\
        );

    \I__4750\ : Span4Mux_v
    port map (
            O => \N__28510\,
            I => \N__28504\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__28507\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__4748\ : Odrv4
    port map (
            O => \N__28504\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__28499\,
            I => \N__28495\
        );

    \I__4746\ : InMux
    port map (
            O => \N__28498\,
            I => \N__28492\
        );

    \I__4745\ : InMux
    port map (
            O => \N__28495\,
            I => \N__28488\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__28492\,
            I => \N__28485\
        );

    \I__4743\ : InMux
    port map (
            O => \N__28491\,
            I => \N__28482\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__28488\,
            I => \N__28477\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__28485\,
            I => \N__28477\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__28482\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__28477\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__28472\,
            I => \N__28468\
        );

    \I__4737\ : InMux
    port map (
            O => \N__28471\,
            I => \N__28465\
        );

    \I__4736\ : InMux
    port map (
            O => \N__28468\,
            I => \N__28460\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__28465\,
            I => \N__28457\
        );

    \I__4734\ : InMux
    port map (
            O => \N__28464\,
            I => \N__28454\
        );

    \I__4733\ : InMux
    port map (
            O => \N__28463\,
            I => \N__28451\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__28460\,
            I => \N__28447\
        );

    \I__4731\ : Span4Mux_v
    port map (
            O => \N__28457\,
            I => \N__28442\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__28454\,
            I => \N__28442\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__28451\,
            I => \N__28439\
        );

    \I__4728\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28436\
        );

    \I__4727\ : Span4Mux_v
    port map (
            O => \N__28447\,
            I => \N__28431\
        );

    \I__4726\ : Span4Mux_h
    port map (
            O => \N__28442\,
            I => \N__28431\
        );

    \I__4725\ : Odrv4
    port map (
            O => \N__28439\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__28436\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4723\ : Odrv4
    port map (
            O => \N__28431\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4722\ : InMux
    port map (
            O => \N__28424\,
            I => \N__28421\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__28421\,
            I => \N__28418\
        );

    \I__4720\ : Span4Mux_v
    port map (
            O => \N__28418\,
            I => \N__28415\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__28415\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\
        );

    \I__4718\ : InMux
    port map (
            O => \N__28412\,
            I => \N__28409\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__28409\,
            I => \N__28406\
        );

    \I__4716\ : Odrv4
    port map (
            O => \N__28406\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\
        );

    \I__4715\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28400\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__28400\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__4713\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28393\
        );

    \I__4712\ : InMux
    port map (
            O => \N__28396\,
            I => \N__28389\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__28393\,
            I => \N__28386\
        );

    \I__4710\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28383\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__28389\,
            I => \N__28380\
        );

    \I__4708\ : Span4Mux_v
    port map (
            O => \N__28386\,
            I => \N__28375\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__28383\,
            I => \N__28375\
        );

    \I__4706\ : Span4Mux_h
    port map (
            O => \N__28380\,
            I => \N__28371\
        );

    \I__4705\ : Span4Mux_h
    port map (
            O => \N__28375\,
            I => \N__28368\
        );

    \I__4704\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28365\
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__28371\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4702\ : Odrv4
    port map (
            O => \N__28368\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__28365\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4700\ : InMux
    port map (
            O => \N__28358\,
            I => \N__28355\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__28355\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__4698\ : CascadeMux
    port map (
            O => \N__28352\,
            I => \N__28348\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__28351\,
            I => \N__28344\
        );

    \I__4696\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28341\
        );

    \I__4695\ : InMux
    port map (
            O => \N__28347\,
            I => \N__28338\
        );

    \I__4694\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28335\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__28341\,
            I => \N__28332\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__28338\,
            I => \N__28327\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__28335\,
            I => \N__28327\
        );

    \I__4690\ : Span4Mux_v
    port map (
            O => \N__28332\,
            I => \N__28323\
        );

    \I__4689\ : Span4Mux_v
    port map (
            O => \N__28327\,
            I => \N__28320\
        );

    \I__4688\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28317\
        );

    \I__4687\ : Odrv4
    port map (
            O => \N__28323\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__28320\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__28317\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4684\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28307\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__28307\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__28304\,
            I => \N__28289\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__28303\,
            I => \N__28286\
        );

    \I__4680\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28274\
        );

    \I__4679\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28274\
        );

    \I__4678\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28269\
        );

    \I__4677\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28269\
        );

    \I__4676\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28266\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28297\,
            I => \N__28255\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28255\
        );

    \I__4673\ : InMux
    port map (
            O => \N__28295\,
            I => \N__28255\
        );

    \I__4672\ : InMux
    port map (
            O => \N__28294\,
            I => \N__28255\
        );

    \I__4671\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28255\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__28292\,
            I => \N__28243\
        );

    \I__4669\ : InMux
    port map (
            O => \N__28289\,
            I => \N__28230\
        );

    \I__4668\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28230\
        );

    \I__4667\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28230\
        );

    \I__4666\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28230\
        );

    \I__4665\ : InMux
    port map (
            O => \N__28283\,
            I => \N__28230\
        );

    \I__4664\ : InMux
    port map (
            O => \N__28282\,
            I => \N__28221\
        );

    \I__4663\ : InMux
    port map (
            O => \N__28281\,
            I => \N__28221\
        );

    \I__4662\ : InMux
    port map (
            O => \N__28280\,
            I => \N__28221\
        );

    \I__4661\ : InMux
    port map (
            O => \N__28279\,
            I => \N__28221\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__28274\,
            I => \N__28216\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__28269\,
            I => \N__28216\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__28266\,
            I => \N__28213\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__28255\,
            I => \N__28210\
        );

    \I__4656\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28205\
        );

    \I__4655\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28205\
        );

    \I__4654\ : InMux
    port map (
            O => \N__28252\,
            I => \N__28196\
        );

    \I__4653\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28196\
        );

    \I__4652\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28196\
        );

    \I__4651\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28196\
        );

    \I__4650\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28183\
        );

    \I__4649\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28183\
        );

    \I__4648\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28183\
        );

    \I__4647\ : InMux
    port map (
            O => \N__28243\,
            I => \N__28183\
        );

    \I__4646\ : InMux
    port map (
            O => \N__28242\,
            I => \N__28183\
        );

    \I__4645\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28183\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__28230\,
            I => \N__28178\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__28221\,
            I => \N__28178\
        );

    \I__4642\ : Span4Mux_h
    port map (
            O => \N__28216\,
            I => \N__28173\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__28213\,
            I => \N__28173\
        );

    \I__4640\ : Span4Mux_v
    port map (
            O => \N__28210\,
            I => \N__28170\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__28205\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__28196\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__28183\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__28178\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__28173\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4634\ : Odrv4
    port map (
            O => \N__28170\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__4633\ : InMux
    port map (
            O => \N__28157\,
            I => \N__28133\
        );

    \I__4632\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28133\
        );

    \I__4631\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28133\
        );

    \I__4630\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28133\
        );

    \I__4629\ : InMux
    port map (
            O => \N__28153\,
            I => \N__28133\
        );

    \I__4628\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28108\
        );

    \I__4627\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28108\
        );

    \I__4626\ : InMux
    port map (
            O => \N__28150\,
            I => \N__28108\
        );

    \I__4625\ : InMux
    port map (
            O => \N__28149\,
            I => \N__28108\
        );

    \I__4624\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28108\
        );

    \I__4623\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28108\
        );

    \I__4622\ : InMux
    port map (
            O => \N__28146\,
            I => \N__28103\
        );

    \I__4621\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28103\
        );

    \I__4620\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28098\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__28133\,
            I => \N__28095\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__28132\,
            I => \N__28091\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__28131\,
            I => \N__28088\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__28130\,
            I => \N__28085\
        );

    \I__4615\ : InMux
    port map (
            O => \N__28129\,
            I => \N__28074\
        );

    \I__4614\ : InMux
    port map (
            O => \N__28128\,
            I => \N__28074\
        );

    \I__4613\ : InMux
    port map (
            O => \N__28127\,
            I => \N__28074\
        );

    \I__4612\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28074\
        );

    \I__4611\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28063\
        );

    \I__4610\ : InMux
    port map (
            O => \N__28124\,
            I => \N__28063\
        );

    \I__4609\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28063\
        );

    \I__4608\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28063\
        );

    \I__4607\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28063\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__28108\,
            I => \N__28058\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__28103\,
            I => \N__28058\
        );

    \I__4604\ : InMux
    port map (
            O => \N__28102\,
            I => \N__28053\
        );

    \I__4603\ : InMux
    port map (
            O => \N__28101\,
            I => \N__28053\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__28098\,
            I => \N__28050\
        );

    \I__4601\ : Span4Mux_v
    port map (
            O => \N__28095\,
            I => \N__28047\
        );

    \I__4600\ : InMux
    port map (
            O => \N__28094\,
            I => \N__28044\
        );

    \I__4599\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28041\
        );

    \I__4598\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28032\
        );

    \I__4597\ : InMux
    port map (
            O => \N__28085\,
            I => \N__28032\
        );

    \I__4596\ : InMux
    port map (
            O => \N__28084\,
            I => \N__28032\
        );

    \I__4595\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28032\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__28074\,
            I => \N__28025\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__28063\,
            I => \N__28025\
        );

    \I__4592\ : Span4Mux_v
    port map (
            O => \N__28058\,
            I => \N__28025\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28018\
        );

    \I__4590\ : Span4Mux_v
    port map (
            O => \N__28050\,
            I => \N__28018\
        );

    \I__4589\ : Span4Mux_v
    port map (
            O => \N__28047\,
            I => \N__28018\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__28044\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__28041\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__28032\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__28025\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__28018\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__4583\ : CascadeMux
    port map (
            O => \N__28007\,
            I => \N__27997\
        );

    \I__4582\ : CascadeMux
    port map (
            O => \N__28006\,
            I => \N__27994\
        );

    \I__4581\ : CascadeMux
    port map (
            O => \N__28005\,
            I => \N__27991\
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__28004\,
            I => \N__27988\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__28003\,
            I => \N__27982\
        );

    \I__4578\ : CascadeMux
    port map (
            O => \N__28002\,
            I => \N__27978\
        );

    \I__4577\ : CascadeMux
    port map (
            O => \N__28001\,
            I => \N__27975\
        );

    \I__4576\ : CascadeMux
    port map (
            O => \N__28000\,
            I => \N__27972\
        );

    \I__4575\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27959\
        );

    \I__4574\ : InMux
    port map (
            O => \N__27994\,
            I => \N__27959\
        );

    \I__4573\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27948\
        );

    \I__4572\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27948\
        );

    \I__4571\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27948\
        );

    \I__4570\ : InMux
    port map (
            O => \N__27986\,
            I => \N__27948\
        );

    \I__4569\ : InMux
    port map (
            O => \N__27985\,
            I => \N__27948\
        );

    \I__4568\ : InMux
    port map (
            O => \N__27982\,
            I => \N__27939\
        );

    \I__4567\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27939\
        );

    \I__4566\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27939\
        );

    \I__4565\ : InMux
    port map (
            O => \N__27975\,
            I => \N__27939\
        );

    \I__4564\ : InMux
    port map (
            O => \N__27972\,
            I => \N__27928\
        );

    \I__4563\ : InMux
    port map (
            O => \N__27971\,
            I => \N__27928\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27970\,
            I => \N__27928\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27969\,
            I => \N__27928\
        );

    \I__4560\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27928\
        );

    \I__4559\ : InMux
    port map (
            O => \N__27967\,
            I => \N__27923\
        );

    \I__4558\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27923\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__27965\,
            I => \N__27919\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__27964\,
            I => \N__27916\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__27959\,
            I => \N__27907\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__27948\,
            I => \N__27907\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__27939\,
            I => \N__27907\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__27928\,
            I => \N__27904\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__27923\,
            I => \N__27900\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27922\,
            I => \N__27895\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27919\,
            I => \N__27895\
        );

    \I__4548\ : InMux
    port map (
            O => \N__27916\,
            I => \N__27890\
        );

    \I__4547\ : InMux
    port map (
            O => \N__27915\,
            I => \N__27890\
        );

    \I__4546\ : CascadeMux
    port map (
            O => \N__27914\,
            I => \N__27887\
        );

    \I__4545\ : Span4Mux_v
    port map (
            O => \N__27907\,
            I => \N__27874\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__27904\,
            I => \N__27874\
        );

    \I__4543\ : InMux
    port map (
            O => \N__27903\,
            I => \N__27871\
        );

    \I__4542\ : Span4Mux_v
    port map (
            O => \N__27900\,
            I => \N__27864\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__27895\,
            I => \N__27864\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__27890\,
            I => \N__27864\
        );

    \I__4539\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27861\
        );

    \I__4538\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27858\
        );

    \I__4537\ : InMux
    port map (
            O => \N__27885\,
            I => \N__27855\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__27884\,
            I => \N__27852\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__27883\,
            I => \N__27849\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__27882\,
            I => \N__27846\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__27881\,
            I => \N__27843\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__27880\,
            I => \N__27840\
        );

    \I__4531\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27837\
        );

    \I__4530\ : Span4Mux_h
    port map (
            O => \N__27874\,
            I => \N__27834\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__27871\,
            I => \N__27831\
        );

    \I__4528\ : Span4Mux_h
    port map (
            O => \N__27864\,
            I => \N__27828\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__27861\,
            I => \N__27825\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27820\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__27855\,
            I => \N__27820\
        );

    \I__4524\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27813\
        );

    \I__4523\ : InMux
    port map (
            O => \N__27849\,
            I => \N__27813\
        );

    \I__4522\ : InMux
    port map (
            O => \N__27846\,
            I => \N__27813\
        );

    \I__4521\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27808\
        );

    \I__4520\ : InMux
    port map (
            O => \N__27840\,
            I => \N__27808\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__27837\,
            I => \N__27805\
        );

    \I__4518\ : Sp12to4
    port map (
            O => \N__27834\,
            I => \N__27802\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__27831\,
            I => \N__27793\
        );

    \I__4516\ : Span4Mux_v
    port map (
            O => \N__27828\,
            I => \N__27793\
        );

    \I__4515\ : Span4Mux_v
    port map (
            O => \N__27825\,
            I => \N__27793\
        );

    \I__4514\ : Span4Mux_v
    port map (
            O => \N__27820\,
            I => \N__27793\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__27813\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__27808\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__27805\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4510\ : Odrv12
    port map (
            O => \N__27802\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__27793\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__4508\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27779\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__27779\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__27776\,
            I => \N__27773\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27769\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27772\,
            I => \N__27766\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__27769\,
            I => \N__27762\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__27766\,
            I => \N__27759\
        );

    \I__4501\ : InMux
    port map (
            O => \N__27765\,
            I => \N__27756\
        );

    \I__4500\ : Span4Mux_h
    port map (
            O => \N__27762\,
            I => \N__27753\
        );

    \I__4499\ : Span4Mux_v
    port map (
            O => \N__27759\,
            I => \N__27748\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__27756\,
            I => \N__27748\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__27753\,
            I => \N__27744\
        );

    \I__4496\ : Span4Mux_h
    port map (
            O => \N__27748\,
            I => \N__27741\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27747\,
            I => \N__27738\
        );

    \I__4494\ : Odrv4
    port map (
            O => \N__27744\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__27741\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__27738\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__27731\,
            I => \N__27728\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27725\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__27725\,
            I => \N__27720\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27717\
        );

    \I__4487\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27713\
        );

    \I__4486\ : Span4Mux_h
    port map (
            O => \N__27720\,
            I => \N__27708\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__27717\,
            I => \N__27708\
        );

    \I__4484\ : InMux
    port map (
            O => \N__27716\,
            I => \N__27704\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__27713\,
            I => \N__27701\
        );

    \I__4482\ : Span4Mux_v
    port map (
            O => \N__27708\,
            I => \N__27698\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27695\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27692\
        );

    \I__4479\ : Span4Mux_h
    port map (
            O => \N__27701\,
            I => \N__27689\
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__27698\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__27695\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4476\ : Odrv4
    port map (
            O => \N__27692\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__27689\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4474\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27677\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__27677\,
            I => \N__27674\
        );

    \I__4472\ : Odrv4
    port map (
            O => \N__27674\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27668\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__27668\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\
        );

    \I__4469\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27661\
        );

    \I__4468\ : InMux
    port map (
            O => \N__27664\,
            I => \N__27658\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__27661\,
            I => \N__27655\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__27658\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__4465\ : Odrv4
    port map (
            O => \N__27655\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__4464\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27646\
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__27649\,
            I => \N__27642\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27646\,
            I => \N__27638\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__27645\,
            I => \N__27635\
        );

    \I__4460\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27630\
        );

    \I__4459\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27630\
        );

    \I__4458\ : Span4Mux_h
    port map (
            O => \N__27638\,
            I => \N__27626\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27623\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__27630\,
            I => \N__27620\
        );

    \I__4455\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27617\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__27626\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__27623\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4452\ : Odrv4
    port map (
            O => \N__27620\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__27617\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__27608\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27602\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__27602\,
            I => \N__27599\
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__27599\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\
        );

    \I__4446\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27593\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__27593\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27590\,
            I => \N__27586\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27589\,
            I => \N__27583\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__27586\,
            I => \N__27580\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__27583\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__4440\ : Odrv12
    port map (
            O => \N__27580\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__4439\ : CascadeMux
    port map (
            O => \N__27575\,
            I => \N__27571\
        );

    \I__4438\ : CascadeMux
    port map (
            O => \N__27574\,
            I => \N__27568\
        );

    \I__4437\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27564\
        );

    \I__4436\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27561\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27557\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__27564\,
            I => \N__27554\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__27561\,
            I => \N__27551\
        );

    \I__4432\ : InMux
    port map (
            O => \N__27560\,
            I => \N__27547\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__27557\,
            I => \N__27544\
        );

    \I__4430\ : Span4Mux_h
    port map (
            O => \N__27554\,
            I => \N__27541\
        );

    \I__4429\ : Span4Mux_v
    port map (
            O => \N__27551\,
            I => \N__27538\
        );

    \I__4428\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27535\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__27547\,
            I => \N__27532\
        );

    \I__4426\ : Span4Mux_v
    port map (
            O => \N__27544\,
            I => \N__27529\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__27541\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__27538\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__27535\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__4422\ : Odrv4
    port map (
            O => \N__27532\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__27529\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27515\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__27515\,
            I => \N__27512\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__27512\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\
        );

    \I__4417\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27506\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__27506\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\
        );

    \I__4415\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27500\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__27500\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27494\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__27494\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\
        );

    \I__4411\ : InMux
    port map (
            O => \N__27491\,
            I => \N__27488\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__27488\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27485\,
            I => \N__27482\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__27482\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__27479\,
            I => \N__27476\
        );

    \I__4406\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27473\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__27473\,
            I => \N__27470\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__27470\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\
        );

    \I__4403\ : InMux
    port map (
            O => \N__27467\,
            I => \N__27464\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__27464\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__27461\,
            I => \N__27458\
        );

    \I__4400\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27454\
        );

    \I__4399\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27450\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27454\,
            I => \N__27447\
        );

    \I__4397\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27444\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__27450\,
            I => \N__27439\
        );

    \I__4395\ : Span4Mux_h
    port map (
            O => \N__27447\,
            I => \N__27436\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__27444\,
            I => \N__27433\
        );

    \I__4393\ : InMux
    port map (
            O => \N__27443\,
            I => \N__27428\
        );

    \I__4392\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27428\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__27439\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__27436\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__27433\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__27428\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4387\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27416\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__27416\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27413\,
            I => \N__27410\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__27410\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\
        );

    \I__4383\ : CascadeMux
    port map (
            O => \N__27407\,
            I => \N__27403\
        );

    \I__4382\ : InMux
    port map (
            O => \N__27406\,
            I => \N__27398\
        );

    \I__4381\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27395\
        );

    \I__4380\ : InMux
    port map (
            O => \N__27402\,
            I => \N__27392\
        );

    \I__4379\ : InMux
    port map (
            O => \N__27401\,
            I => \N__27388\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__27398\,
            I => \N__27385\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__27395\,
            I => \N__27382\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__27392\,
            I => \N__27379\
        );

    \I__4375\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27376\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__27388\,
            I => \N__27373\
        );

    \I__4373\ : Span4Mux_h
    port map (
            O => \N__27385\,
            I => \N__27370\
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__27382\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__27379\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__27376\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4369\ : Odrv12
    port map (
            O => \N__27373\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4368\ : Odrv4
    port map (
            O => \N__27370\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4367\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27356\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__27356\,
            I => \N__27353\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__27353\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\
        );

    \I__4364\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27347\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__27347\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\
        );

    \I__4362\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27341\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__27341\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\
        );

    \I__4360\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27335\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__27335\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\
        );

    \I__4358\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27329\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__27329\,
            I => \N__27326\
        );

    \I__4356\ : Odrv12
    port map (
            O => \N__27326\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_10\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__27323\,
            I => \N__27320\
        );

    \I__4354\ : InMux
    port map (
            O => \N__27320\,
            I => \N__27317\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__27317\,
            I => \N__27314\
        );

    \I__4352\ : Odrv4
    port map (
            O => \N__27314\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\
        );

    \I__4351\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27308\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__27308\,
            I => \N__27305\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__27305\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__4348\ : InMux
    port map (
            O => \N__27302\,
            I => \N__27298\
        );

    \I__4347\ : InMux
    port map (
            O => \N__27301\,
            I => \N__27294\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__27298\,
            I => \N__27290\
        );

    \I__4345\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27287\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__27294\,
            I => \N__27284\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__27293\,
            I => \N__27281\
        );

    \I__4342\ : Span4Mux_v
    port map (
            O => \N__27290\,
            I => \N__27276\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__27287\,
            I => \N__27276\
        );

    \I__4340\ : Span4Mux_h
    port map (
            O => \N__27284\,
            I => \N__27272\
        );

    \I__4339\ : InMux
    port map (
            O => \N__27281\,
            I => \N__27269\
        );

    \I__4338\ : Span4Mux_h
    port map (
            O => \N__27276\,
            I => \N__27266\
        );

    \I__4337\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27263\
        );

    \I__4336\ : Span4Mux_v
    port map (
            O => \N__27272\,
            I => \N__27260\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__27269\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__27266\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__27263\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__27260\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4331\ : InMux
    port map (
            O => \N__27251\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\
        );

    \I__4330\ : InMux
    port map (
            O => \N__27248\,
            I => \bfn_11_11_0_\
        );

    \I__4329\ : InMux
    port map (
            O => \N__27245\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\
        );

    \I__4328\ : InMux
    port map (
            O => \N__27242\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\
        );

    \I__4327\ : InMux
    port map (
            O => \N__27239\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\
        );

    \I__4326\ : InMux
    port map (
            O => \N__27236\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\
        );

    \I__4325\ : InMux
    port map (
            O => \N__27233\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\
        );

    \I__4324\ : InMux
    port map (
            O => \N__27230\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\
        );

    \I__4323\ : InMux
    port map (
            O => \N__27227\,
            I => \N__27223\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__27226\,
            I => \N__27220\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__27223\,
            I => \N__27215\
        );

    \I__4320\ : InMux
    port map (
            O => \N__27220\,
            I => \N__27212\
        );

    \I__4319\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27209\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__27218\,
            I => \N__27205\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__27215\,
            I => \N__27200\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__27212\,
            I => \N__27200\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__27209\,
            I => \N__27197\
        );

    \I__4314\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27192\
        );

    \I__4313\ : InMux
    port map (
            O => \N__27205\,
            I => \N__27192\
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__27200\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__4311\ : Odrv4
    port map (
            O => \N__27197\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__27192\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__4309\ : InMux
    port map (
            O => \N__27185\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_31\
        );

    \I__4308\ : InMux
    port map (
            O => \N__27182\,
            I => \N__27179\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__27179\,
            I => \N__27176\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__27176\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\
        );

    \I__4305\ : InMux
    port map (
            O => \N__27173\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\
        );

    \I__4304\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27167\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__27167\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\
        );

    \I__4302\ : InMux
    port map (
            O => \N__27164\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\
        );

    \I__4301\ : InMux
    port map (
            O => \N__27161\,
            I => \bfn_11_10_0_\
        );

    \I__4300\ : InMux
    port map (
            O => \N__27158\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\
        );

    \I__4299\ : InMux
    port map (
            O => \N__27155\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\
        );

    \I__4298\ : InMux
    port map (
            O => \N__27152\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\
        );

    \I__4297\ : InMux
    port map (
            O => \N__27149\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\
        );

    \I__4296\ : InMux
    port map (
            O => \N__27146\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\
        );

    \I__4295\ : InMux
    port map (
            O => \N__27143\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\
        );

    \I__4294\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27137\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__27137\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_6\
        );

    \I__4292\ : InMux
    port map (
            O => \N__27134\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\
        );

    \I__4291\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27128\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__27128\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_7\
        );

    \I__4289\ : InMux
    port map (
            O => \N__27125\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\
        );

    \I__4288\ : InMux
    port map (
            O => \N__27122\,
            I => \N__27119\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__27119\,
            I => \N__27116\
        );

    \I__4286\ : Odrv12
    port map (
            O => \N__27116\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\
        );

    \I__4285\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27110\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__27110\,
            I => \N__27107\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__27107\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_8\
        );

    \I__4282\ : InMux
    port map (
            O => \N__27104\,
            I => \bfn_11_9_0_\
        );

    \I__4281\ : InMux
    port map (
            O => \N__27101\,
            I => \N__27098\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__27095\
        );

    \I__4279\ : Odrv12
    port map (
            O => \N__27095\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\
        );

    \I__4278\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27089\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__27089\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_9\
        );

    \I__4276\ : InMux
    port map (
            O => \N__27086\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\
        );

    \I__4275\ : InMux
    port map (
            O => \N__27083\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\
        );

    \I__4274\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27077\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__27077\,
            I => \N__27074\
        );

    \I__4272\ : Span4Mux_v
    port map (
            O => \N__27074\,
            I => \N__27071\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__27071\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_11\
        );

    \I__4270\ : InMux
    port map (
            O => \N__27068\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\
        );

    \I__4269\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27062\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__27062\,
            I => \N__27059\
        );

    \I__4267\ : Odrv4
    port map (
            O => \N__27059\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\
        );

    \I__4266\ : InMux
    port map (
            O => \N__27056\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\
        );

    \I__4265\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27050\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__27050\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27047\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\
        );

    \I__4262\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27041\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__27041\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\
        );

    \I__4260\ : InMux
    port map (
            O => \N__27038\,
            I => \N__27035\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__27035\,
            I => \N__27032\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__27032\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__27029\,
            I => \N__27026\
        );

    \I__4256\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27023\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__27023\,
            I => \N__27020\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__27020\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__4253\ : InMux
    port map (
            O => \N__27017\,
            I => \N__27014\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__27014\,
            I => \N__27011\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__27011\,
            I => \N__27007\
        );

    \I__4250\ : InMux
    port map (
            O => \N__27010\,
            I => \N__27004\
        );

    \I__4249\ : Odrv4
    port map (
            O => \N__27007\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__27004\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__4247\ : InMux
    port map (
            O => \N__26999\,
            I => \N__26996\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__26996\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\
        );

    \I__4245\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26990\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__26990\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\
        );

    \I__4243\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26984\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__26984\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\
        );

    \I__4241\ : InMux
    port map (
            O => \N__26981\,
            I => \N__26978\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__26978\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\
        );

    \I__4239\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26972\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__26972\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_4\
        );

    \I__4237\ : InMux
    port map (
            O => \N__26969\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\
        );

    \I__4236\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26963\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__26963\,
            I => \N__26960\
        );

    \I__4234\ : Odrv4
    port map (
            O => \N__26960\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_5\
        );

    \I__4233\ : InMux
    port map (
            O => \N__26957\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__26954\,
            I => \N__26951\
        );

    \I__4231\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26948\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__26948\,
            I => \N__26945\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__26945\,
            I => \N__26942\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__26942\,
            I => \current_shift_inst.PI_CTRL.integrator_i_21\
        );

    \I__4227\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26901\
        );

    \I__4226\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26901\
        );

    \I__4225\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26901\
        );

    \I__4224\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26901\
        );

    \I__4223\ : InMux
    port map (
            O => \N__26935\,
            I => \N__26892\
        );

    \I__4222\ : InMux
    port map (
            O => \N__26934\,
            I => \N__26892\
        );

    \I__4221\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26892\
        );

    \I__4220\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26892\
        );

    \I__4219\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26883\
        );

    \I__4218\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26883\
        );

    \I__4217\ : InMux
    port map (
            O => \N__26929\,
            I => \N__26883\
        );

    \I__4216\ : InMux
    port map (
            O => \N__26928\,
            I => \N__26883\
        );

    \I__4215\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26874\
        );

    \I__4214\ : InMux
    port map (
            O => \N__26926\,
            I => \N__26874\
        );

    \I__4213\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26874\
        );

    \I__4212\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26874\
        );

    \I__4211\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26869\
        );

    \I__4210\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26869\
        );

    \I__4209\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26860\
        );

    \I__4208\ : InMux
    port map (
            O => \N__26920\,
            I => \N__26860\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26860\
        );

    \I__4206\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26860\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26851\
        );

    \I__4204\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26851\
        );

    \I__4203\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26851\
        );

    \I__4202\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26851\
        );

    \I__4201\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26842\
        );

    \I__4200\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26842\
        );

    \I__4199\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26842\
        );

    \I__4198\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26842\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__26901\,
            I => \N__26839\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__26892\,
            I => \N__26836\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__26883\,
            I => \N__26831\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__26874\,
            I => \N__26831\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__26869\,
            I => \N__26828\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__26860\,
            I => \N__26825\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__26851\,
            I => \N__26820\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__26842\,
            I => \N__26820\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__26839\,
            I => \N__26817\
        );

    \I__4188\ : Span4Mux_h
    port map (
            O => \N__26836\,
            I => \N__26814\
        );

    \I__4187\ : Span4Mux_h
    port map (
            O => \N__26831\,
            I => \N__26811\
        );

    \I__4186\ : Span4Mux_v
    port map (
            O => \N__26828\,
            I => \N__26806\
        );

    \I__4185\ : Span4Mux_v
    port map (
            O => \N__26825\,
            I => \N__26806\
        );

    \I__4184\ : Span4Mux_h
    port map (
            O => \N__26820\,
            I => \N__26803\
        );

    \I__4183\ : Span4Mux_v
    port map (
            O => \N__26817\,
            I => \N__26798\
        );

    \I__4182\ : Span4Mux_v
    port map (
            O => \N__26814\,
            I => \N__26798\
        );

    \I__4181\ : Span4Mux_v
    port map (
            O => \N__26811\,
            I => \N__26795\
        );

    \I__4180\ : Odrv4
    port map (
            O => \N__26806\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4179\ : Odrv4
    port map (
            O => \N__26803\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4178\ : Odrv4
    port map (
            O => \N__26798\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4177\ : Odrv4
    port map (
            O => \N__26795\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4176\ : InMux
    port map (
            O => \N__26786\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__26783\,
            I => \N__26780\
        );

    \I__4174\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26776\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26779\,
            I => \N__26773\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__26776\,
            I => \N__26770\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__26773\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__4170\ : Odrv4
    port map (
            O => \N__26770\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26759\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26756\
        );

    \I__4167\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26751\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26751\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__26759\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__26756\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__26751\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__26744\,
            I => \delay_measurement_inst.N_39_cascade_\
        );

    \I__4161\ : InMux
    port map (
            O => \N__26741\,
            I => \N__26738\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__26738\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4159\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26732\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__26732\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__26729\,
            I => \N__26726\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26723\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26723\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_26\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26717\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__26717\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26714\,
            I => \N__26711\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26711\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26705\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__26705\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__4148\ : InMux
    port map (
            O => \N__26702\,
            I => \N__26699\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__26699\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2\
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__26696\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_\
        );

    \I__4145\ : InMux
    port map (
            O => \N__26693\,
            I => \N__26690\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__26690\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26687\,
            I => \N__26684\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__26684\,
            I => \N__26681\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__26681\,
            I => \N__26677\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26674\
        );

    \I__4139\ : Odrv4
    port map (
            O => \N__26677\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26674\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__4137\ : InMux
    port map (
            O => \N__26669\,
            I => \N__26665\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26662\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__26665\,
            I => \delay_measurement_inst.elapsed_time_hc_27\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26662\,
            I => \delay_measurement_inst.elapsed_time_hc_27\
        );

    \I__4133\ : IoInMux
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__26654\,
            I => \N__26651\
        );

    \I__4131\ : Span4Mux_s3_v
    port map (
            O => \N__26651\,
            I => \N__26648\
        );

    \I__4130\ : Sp12to4
    port map (
            O => \N__26648\,
            I => \N__26645\
        );

    \I__4129\ : Odrv12
    port map (
            O => \N__26645\,
            I => s3_phy_c
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__26642\,
            I => \N__26638\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__26641\,
            I => \N__26635\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26629\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26635\,
            I => \N__26629\
        );

    \I__4124\ : InMux
    port map (
            O => \N__26634\,
            I => \N__26626\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26629\,
            I => \N__26623\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__26626\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__26623\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__4120\ : InMux
    port map (
            O => \N__26618\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__26615\,
            I => \N__26612\
        );

    \I__4118\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26608\
        );

    \I__4117\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26604\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__26608\,
            I => \N__26601\
        );

    \I__4115\ : InMux
    port map (
            O => \N__26607\,
            I => \N__26598\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__26604\,
            I => \N__26593\
        );

    \I__4113\ : Span4Mux_h
    port map (
            O => \N__26601\,
            I => \N__26593\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__26598\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__26593\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26588\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26579\
        );

    \I__4108\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26579\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__26579\,
            I => \N__26575\
        );

    \I__4106\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26572\
        );

    \I__4105\ : Span4Mux_h
    port map (
            O => \N__26575\,
            I => \N__26569\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__26572\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__26569\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__4102\ : InMux
    port map (
            O => \N__26564\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__4101\ : CascadeMux
    port map (
            O => \N__26561\,
            I => \N__26558\
        );

    \I__4100\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26554\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__26557\,
            I => \N__26550\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__26554\,
            I => \N__26547\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26544\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26541\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__26547\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__26544\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__26541\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4092\ : InMux
    port map (
            O => \N__26534\,
            I => \bfn_10_20_0_\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__26531\,
            I => \N__26528\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26525\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__26525\,
            I => \N__26520\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__26524\,
            I => \N__26517\
        );

    \I__4087\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26514\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__26520\,
            I => \N__26511\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26508\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__26514\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__26511\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__26508\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4081\ : InMux
    port map (
            O => \N__26501\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__4079\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26491\
        );

    \I__4078\ : InMux
    port map (
            O => \N__26494\,
            I => \N__26488\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__26491\,
            I => \N__26482\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__26488\,
            I => \N__26482\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26487\,
            I => \N__26479\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__26482\,
            I => \N__26476\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26479\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__26476\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__4071\ : InMux
    port map (
            O => \N__26471\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__4070\ : InMux
    port map (
            O => \N__26468\,
            I => \N__26461\
        );

    \I__4069\ : InMux
    port map (
            O => \N__26467\,
            I => \N__26461\
        );

    \I__4068\ : InMux
    port map (
            O => \N__26466\,
            I => \N__26458\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__26461\,
            I => \N__26455\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__26458\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__4065\ : Odrv4
    port map (
            O => \N__26455\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__4064\ : InMux
    port map (
            O => \N__26450\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__4063\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26443\
        );

    \I__4062\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26440\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__26443\,
            I => \N__26437\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__26440\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__4059\ : Odrv4
    port map (
            O => \N__26437\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26432\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__4057\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26422\
        );

    \I__4056\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26422\
        );

    \I__4055\ : InMux
    port map (
            O => \N__26427\,
            I => \N__26419\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__26422\,
            I => \N__26416\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26419\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__26416\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4051\ : InMux
    port map (
            O => \N__26411\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__4050\ : CascadeMux
    port map (
            O => \N__26408\,
            I => \N__26404\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__26407\,
            I => \N__26401\
        );

    \I__4048\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26395\
        );

    \I__4047\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26395\
        );

    \I__4046\ : InMux
    port map (
            O => \N__26400\,
            I => \N__26392\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__26395\,
            I => \N__26389\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__26392\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__26389\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4042\ : InMux
    port map (
            O => \N__26384\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__26381\,
            I => \N__26378\
        );

    \I__4040\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26374\
        );

    \I__4039\ : InMux
    port map (
            O => \N__26377\,
            I => \N__26370\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__26374\,
            I => \N__26367\
        );

    \I__4037\ : InMux
    port map (
            O => \N__26373\,
            I => \N__26364\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__26370\,
            I => \N__26359\
        );

    \I__4035\ : Span4Mux_h
    port map (
            O => \N__26367\,
            I => \N__26359\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__26364\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__26359\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4032\ : InMux
    port map (
            O => \N__26354\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__4031\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26345\
        );

    \I__4030\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26345\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__26345\,
            I => \N__26341\
        );

    \I__4028\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26338\
        );

    \I__4027\ : Span4Mux_h
    port map (
            O => \N__26341\,
            I => \N__26335\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__26338\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__26335\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4024\ : InMux
    port map (
            O => \N__26330\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__4023\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26323\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__26326\,
            I => \N__26319\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__26323\,
            I => \N__26316\
        );

    \I__4020\ : InMux
    port map (
            O => \N__26322\,
            I => \N__26313\
        );

    \I__4019\ : InMux
    port map (
            O => \N__26319\,
            I => \N__26310\
        );

    \I__4018\ : Span4Mux_h
    port map (
            O => \N__26316\,
            I => \N__26307\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__26313\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__26310\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4015\ : Odrv4
    port map (
            O => \N__26307\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4014\ : InMux
    port map (
            O => \N__26300\,
            I => \bfn_10_19_0_\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__26297\,
            I => \N__26294\
        );

    \I__4012\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__26291\,
            I => \N__26286\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__26290\,
            I => \N__26283\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26280\
        );

    \I__4008\ : Span4Mux_h
    port map (
            O => \N__26286\,
            I => \N__26277\
        );

    \I__4007\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26274\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__26280\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4005\ : Odrv4
    port map (
            O => \N__26277\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__26274\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4003\ : InMux
    port map (
            O => \N__26267\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__26264\,
            I => \N__26260\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__26263\,
            I => \N__26257\
        );

    \I__4000\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26251\
        );

    \I__3999\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26251\
        );

    \I__3998\ : InMux
    port map (
            O => \N__26256\,
            I => \N__26248\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__26251\,
            I => \N__26245\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__26248\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__26245\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__3994\ : InMux
    port map (
            O => \N__26240\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__3993\ : InMux
    port map (
            O => \N__26237\,
            I => \N__26230\
        );

    \I__3992\ : InMux
    port map (
            O => \N__26236\,
            I => \N__26230\
        );

    \I__3991\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26227\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__26230\,
            I => \N__26224\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__26227\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__3988\ : Odrv4
    port map (
            O => \N__26224\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__3987\ : InMux
    port map (
            O => \N__26219\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__3986\ : InMux
    port map (
            O => \N__26216\,
            I => \N__26209\
        );

    \I__3985\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26209\
        );

    \I__3984\ : InMux
    port map (
            O => \N__26214\,
            I => \N__26206\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__26209\,
            I => \N__26203\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__26206\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__26203\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__3980\ : InMux
    port map (
            O => \N__26198\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__26195\,
            I => \N__26191\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__26194\,
            I => \N__26188\
        );

    \I__3977\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26183\
        );

    \I__3976\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26183\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26179\
        );

    \I__3974\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26176\
        );

    \I__3973\ : Span4Mux_h
    port map (
            O => \N__26179\,
            I => \N__26173\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__26176\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__3971\ : Odrv4
    port map (
            O => \N__26173\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__3970\ : InMux
    port map (
            O => \N__26168\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__3969\ : CascadeMux
    port map (
            O => \N__26165\,
            I => \N__26161\
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__26164\,
            I => \N__26158\
        );

    \I__3967\ : InMux
    port map (
            O => \N__26161\,
            I => \N__26152\
        );

    \I__3966\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26152\
        );

    \I__3965\ : InMux
    port map (
            O => \N__26157\,
            I => \N__26149\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__26152\,
            I => \N__26146\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__26149\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__26146\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__3961\ : InMux
    port map (
            O => \N__26141\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__3960\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26131\
        );

    \I__3959\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26131\
        );

    \I__3958\ : InMux
    port map (
            O => \N__26136\,
            I => \N__26128\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__26131\,
            I => \N__26125\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__26128\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__26125\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__3954\ : InMux
    port map (
            O => \N__26120\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__3953\ : InMux
    port map (
            O => \N__26117\,
            I => \N__26111\
        );

    \I__3952\ : InMux
    port map (
            O => \N__26116\,
            I => \N__26111\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__26111\,
            I => \N__26107\
        );

    \I__3950\ : InMux
    port map (
            O => \N__26110\,
            I => \N__26104\
        );

    \I__3949\ : Span4Mux_h
    port map (
            O => \N__26107\,
            I => \N__26101\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__26104\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__26101\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__3946\ : InMux
    port map (
            O => \N__26096\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__3945\ : InMux
    port map (
            O => \N__26093\,
            I => \N__26090\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__26090\,
            I => \N__26086\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__26089\,
            I => \N__26082\
        );

    \I__3942\ : Span4Mux_v
    port map (
            O => \N__26086\,
            I => \N__26079\
        );

    \I__3941\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26076\
        );

    \I__3940\ : InMux
    port map (
            O => \N__26082\,
            I => \N__26073\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__26079\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__26076\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__26073\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__3936\ : InMux
    port map (
            O => \N__26066\,
            I => \bfn_10_18_0_\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__26063\,
            I => \N__26060\
        );

    \I__3934\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26057\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__26057\,
            I => \N__26052\
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__26056\,
            I => \N__26049\
        );

    \I__3931\ : InMux
    port map (
            O => \N__26055\,
            I => \N__26046\
        );

    \I__3930\ : Span4Mux_h
    port map (
            O => \N__26052\,
            I => \N__26043\
        );

    \I__3929\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26040\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__26046\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__26043\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__26040\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__3925\ : InMux
    port map (
            O => \N__26033\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__3924\ : CascadeMux
    port map (
            O => \N__26030\,
            I => \N__26026\
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__26029\,
            I => \N__26023\
        );

    \I__3922\ : InMux
    port map (
            O => \N__26026\,
            I => \N__26017\
        );

    \I__3921\ : InMux
    port map (
            O => \N__26023\,
            I => \N__26017\
        );

    \I__3920\ : InMux
    port map (
            O => \N__26022\,
            I => \N__26014\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__26017\,
            I => \N__26011\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__26014\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__26011\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__3916\ : InMux
    port map (
            O => \N__26006\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__3915\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25996\
        );

    \I__3914\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25996\
        );

    \I__3913\ : InMux
    port map (
            O => \N__26001\,
            I => \N__25993\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__25996\,
            I => \N__25990\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__25993\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__25990\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25985\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__25982\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_\
        );

    \I__3907\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25975\
        );

    \I__3906\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25971\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__25975\,
            I => \N__25968\
        );

    \I__3904\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25965\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__25971\,
            I => \N__25960\
        );

    \I__3902\ : Span4Mux_v
    port map (
            O => \N__25968\,
            I => \N__25960\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__25965\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__25960\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25952\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__25952\,
            I => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__25949\,
            I => \phase_controller_inst1.stoper_hc.time_passed11_cascade_\
        );

    \I__3896\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25943\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__25943\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__3894\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25936\
        );

    \I__3893\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25933\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__25936\,
            I => \N__25930\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__25933\,
            I => \N__25925\
        );

    \I__3890\ : Span4Mux_h
    port map (
            O => \N__25930\,
            I => \N__25925\
        );

    \I__3889\ : Odrv4
    port map (
            O => \N__25925\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3888\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25918\
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__25921\,
            I => \N__25915\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__25918\,
            I => \N__25912\
        );

    \I__3885\ : InMux
    port map (
            O => \N__25915\,
            I => \N__25909\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__25912\,
            I => \N__25905\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__25909\,
            I => \N__25902\
        );

    \I__3882\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25899\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__25905\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__25902\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__25899\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__3878\ : InMux
    port map (
            O => \N__25892\,
            I => \bfn_10_17_0_\
        );

    \I__3877\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25886\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__25886\,
            I => \N__25883\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__25883\,
            I => \N__25879\
        );

    \I__3874\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25876\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__25879\,
            I => \N__25872\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__25876\,
            I => \N__25869\
        );

    \I__3871\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25866\
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__25872\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__25869\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__25866\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__3867\ : InMux
    port map (
            O => \N__25859\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__3866\ : InMux
    port map (
            O => \N__25856\,
            I => \N__25849\
        );

    \I__3865\ : InMux
    port map (
            O => \N__25855\,
            I => \N__25849\
        );

    \I__3864\ : InMux
    port map (
            O => \N__25854\,
            I => \N__25846\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__25849\,
            I => \N__25843\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__25846\,
            I => \N__25838\
        );

    \I__3861\ : Span4Mux_v
    port map (
            O => \N__25843\,
            I => \N__25838\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__25838\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__3859\ : InMux
    port map (
            O => \N__25835\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__25832\,
            I => \N__25829\
        );

    \I__3857\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25825\
        );

    \I__3856\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25821\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__25825\,
            I => \N__25818\
        );

    \I__3854\ : InMux
    port map (
            O => \N__25824\,
            I => \N__25815\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__25821\,
            I => \N__25812\
        );

    \I__3852\ : Span4Mux_v
    port map (
            O => \N__25818\,
            I => \N__25809\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__25815\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__25812\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__25809\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__3848\ : InMux
    port map (
            O => \N__25802\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__25799\,
            I => \N__25796\
        );

    \I__3846\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__25793\,
            I => \current_shift_inst.PI_CTRL.integrator_i_23\
        );

    \I__3844\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25787\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__25787\,
            I => \current_shift_inst.PI_CTRL.integrator_i_28\
        );

    \I__3842\ : InMux
    port map (
            O => \N__25784\,
            I => \N__25781\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__25781\,
            I => \current_shift_inst.PI_CTRL.integrator_i_30\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__25778\,
            I => \N__25775\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__25772\,
            I => \current_shift_inst.PI_CTRL.integrator_i_29\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25769\,
            I => \N__25766\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__25766\,
            I => \N__25763\
        );

    \I__3835\ : Odrv12
    port map (
            O => \N__25763\,
            I => \current_shift_inst.PI_CTRL.integrator_i_6\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__25760\,
            I => \N__25757\
        );

    \I__3833\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__25754\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\
        );

    \I__3831\ : InMux
    port map (
            O => \N__25751\,
            I => \bfn_10_13_0_\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__3829\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25742\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__25742\,
            I => \N__25739\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__25739\,
            I => \N__25736\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__25736\,
            I => \N__25733\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__25733\,
            I => \current_shift_inst.PI_CTRL.integrator_i_24\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25727\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__25727\,
            I => \N__25724\
        );

    \I__3822\ : Odrv4
    port map (
            O => \N__25724\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__3821\ : InMux
    port map (
            O => \N__25721\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__25718\,
            I => \N__25715\
        );

    \I__3819\ : InMux
    port map (
            O => \N__25715\,
            I => \N__25712\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__25712\,
            I => \N__25709\
        );

    \I__3817\ : Span4Mux_v
    port map (
            O => \N__25709\,
            I => \N__25706\
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__25706\,
            I => \current_shift_inst.PI_CTRL.integrator_i_25\
        );

    \I__3815\ : InMux
    port map (
            O => \N__25703\,
            I => \N__25700\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__25700\,
            I => \N__25697\
        );

    \I__3813\ : Span4Mux_h
    port map (
            O => \N__25697\,
            I => \N__25694\
        );

    \I__3812\ : Odrv4
    port map (
            O => \N__25694\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__3811\ : InMux
    port map (
            O => \N__25691\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__25688\,
            I => \N__25685\
        );

    \I__3809\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25682\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__25682\,
            I => \current_shift_inst.PI_CTRL.integrator_i_26\
        );

    \I__3807\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25676\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__25676\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__3805\ : InMux
    port map (
            O => \N__25673\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__25670\,
            I => \N__25667\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25667\,
            I => \N__25664\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__25664\,
            I => \current_shift_inst.PI_CTRL.integrator_i_27\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25658\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__25658\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25655\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25652\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\
        );

    \I__3797\ : InMux
    port map (
            O => \N__25649\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25646\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25643\,
            I => \bfn_10_14_0_\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__25640\,
            I => \N__25637\
        );

    \I__3793\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25634\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__25634\,
            I => \N__25631\
        );

    \I__3791\ : Odrv4
    port map (
            O => \N__25631\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__3790\ : InMux
    port map (
            O => \N__25628\,
            I => \bfn_10_12_0_\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__25625\,
            I => \N__25622\
        );

    \I__3788\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25619\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__25619\,
            I => \N__25616\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__25616\,
            I => \N__25613\
        );

    \I__3785\ : Span4Mux_h
    port map (
            O => \N__25613\,
            I => \N__25610\
        );

    \I__3784\ : Odrv4
    port map (
            O => \N__25610\,
            I => \current_shift_inst.PI_CTRL.integrator_i_16\
        );

    \I__3783\ : InMux
    port map (
            O => \N__25607\,
            I => \N__25604\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__25604\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__3781\ : InMux
    port map (
            O => \N__25601\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__25598\,
            I => \N__25595\
        );

    \I__3779\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25592\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__25589\,
            I => \N__25586\
        );

    \I__3776\ : Span4Mux_h
    port map (
            O => \N__25586\,
            I => \N__25583\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__25583\,
            I => \current_shift_inst.PI_CTRL.integrator_i_17\
        );

    \I__3774\ : CascadeMux
    port map (
            O => \N__25580\,
            I => \N__25577\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25577\,
            I => \N__25574\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__25574\,
            I => \N__25571\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__25571\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__3770\ : InMux
    port map (
            O => \N__25568\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__25565\,
            I => \N__25562\
        );

    \I__3768\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25559\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__25559\,
            I => \N__25556\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__25556\,
            I => \N__25553\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__25553\,
            I => \current_shift_inst.PI_CTRL.integrator_i_18\
        );

    \I__3764\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25547\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__25547\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25544\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__25541\,
            I => \N__25538\
        );

    \I__3760\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25535\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__25535\,
            I => \N__25532\
        );

    \I__3758\ : Span4Mux_h
    port map (
            O => \N__25532\,
            I => \N__25529\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__25529\,
            I => \current_shift_inst.PI_CTRL.integrator_i_19\
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__25526\,
            I => \N__25523\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__25520\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25517\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__25514\,
            I => \N__25511\
        );

    \I__3751\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25508\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__25508\,
            I => \N__25505\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__25505\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25502\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25496\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__25496\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__3745\ : InMux
    port map (
            O => \N__25493\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__25490\,
            I => \N__25487\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25487\,
            I => \N__25484\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__25484\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25481\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\
        );

    \I__3740\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25475\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__25475\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__3738\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25469\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__25469\,
            I => \N__25466\
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__25466\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__25463\,
            I => \N__25460\
        );

    \I__3734\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25457\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__25457\,
            I => \N__25454\
        );

    \I__3732\ : Span4Mux_v
    port map (
            O => \N__25454\,
            I => \N__25451\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__25451\,
            I => \current_shift_inst.PI_CTRL.integrator_i_8\
        );

    \I__3730\ : InMux
    port map (
            O => \N__25448\,
            I => \N__25445\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__25445\,
            I => \N__25442\
        );

    \I__3728\ : Span4Mux_h
    port map (
            O => \N__25442\,
            I => \N__25439\
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__25439\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__3726\ : InMux
    port map (
            O => \N__25436\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\
        );

    \I__3725\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25430\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__25430\,
            I => \N__25427\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__25427\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__25424\,
            I => \N__25421\
        );

    \I__3721\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25418\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25418\,
            I => \N__25415\
        );

    \I__3719\ : Span4Mux_v
    port map (
            O => \N__25415\,
            I => \N__25412\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__25412\,
            I => \current_shift_inst.PI_CTRL.integrator_i_9\
        );

    \I__3717\ : InMux
    port map (
            O => \N__25409\,
            I => \N__25406\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__25406\,
            I => \N__25403\
        );

    \I__3715\ : Span4Mux_h
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__25400\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__3713\ : InMux
    port map (
            O => \N__25397\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\
        );

    \I__3712\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__25391\,
            I => \N__25388\
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__25388\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__25385\,
            I => \N__25382\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25379\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__3706\ : Span4Mux_v
    port map (
            O => \N__25376\,
            I => \N__25373\
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__25373\,
            I => \current_shift_inst.PI_CTRL.integrator_i_10\
        );

    \I__3704\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25367\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__25367\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__3702\ : InMux
    port map (
            O => \N__25364\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\
        );

    \I__3701\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25358\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__25358\,
            I => \N__25355\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__25355\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\
        );

    \I__3698\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25349\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__25349\,
            I => \N__25346\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__25346\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__3695\ : InMux
    port map (
            O => \N__25343\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__25340\,
            I => \N__25337\
        );

    \I__3693\ : InMux
    port map (
            O => \N__25337\,
            I => \N__25334\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__25334\,
            I => \N__25331\
        );

    \I__3691\ : Span4Mux_h
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__3690\ : Odrv4
    port map (
            O => \N__25328\,
            I => \current_shift_inst.PI_CTRL.integrator_i_12\
        );

    \I__3689\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25322\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25319\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__25319\,
            I => \N__25316\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__25316\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__3685\ : InMux
    port map (
            O => \N__25313\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__25310\,
            I => \N__25307\
        );

    \I__3683\ : InMux
    port map (
            O => \N__25307\,
            I => \N__25304\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__25304\,
            I => \N__25301\
        );

    \I__3681\ : Span4Mux_v
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__25298\,
            I => \current_shift_inst.PI_CTRL.integrator_i_13\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__25295\,
            I => \N__25292\
        );

    \I__3678\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25289\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__25289\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__3676\ : InMux
    port map (
            O => \N__25286\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\
        );

    \I__3675\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25280\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__25280\,
            I => \N__25277\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__25277\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__3672\ : InMux
    port map (
            O => \N__25274\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__25271\,
            I => \N__25268\
        );

    \I__3670\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25265\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__25265\,
            I => \N__25262\
        );

    \I__3668\ : Span4Mux_h
    port map (
            O => \N__25262\,
            I => \N__25259\
        );

    \I__3667\ : Odrv4
    port map (
            O => \N__25259\,
            I => \current_shift_inst.PI_CTRL.integrator_i_15\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__25256\,
            I => \N__25253\
        );

    \I__3665\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25249\
        );

    \I__3664\ : InMux
    port map (
            O => \N__25252\,
            I => \N__25246\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__25249\,
            I => \N__25241\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__25246\,
            I => \N__25241\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__25241\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__3660\ : CascadeMux
    port map (
            O => \N__25238\,
            I => \N__25235\
        );

    \I__3659\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25232\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__25232\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\
        );

    \I__3657\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25226\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__25226\,
            I => \N__25223\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__25223\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\
        );

    \I__3654\ : InMux
    port map (
            O => \N__25220\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\
        );

    \I__3653\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25214\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__25214\,
            I => \N__25211\
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__25211\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__25208\,
            I => \N__25205\
        );

    \I__3649\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25202\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__25202\,
            I => \N__25199\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__25199\,
            I => \current_shift_inst.PI_CTRL.integrator_i_1\
        );

    \I__3646\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25193\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__25193\,
            I => \N__25190\
        );

    \I__3644\ : Span4Mux_v
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__25187\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\
        );

    \I__3642\ : InMux
    port map (
            O => \N__25184\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\
        );

    \I__3641\ : InMux
    port map (
            O => \N__25181\,
            I => \N__25178\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__25178\,
            I => \N__25175\
        );

    \I__3639\ : Odrv4
    port map (
            O => \N__25175\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__25172\,
            I => \N__25169\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25166\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__25166\,
            I => \N__25163\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__25163\,
            I => \current_shift_inst.PI_CTRL.integrator_i_2\
        );

    \I__3634\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25157\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__25157\,
            I => \N__25154\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__25154\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__3631\ : InMux
    port map (
            O => \N__25151\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\
        );

    \I__3630\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25145\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__25145\,
            I => \N__25142\
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__25142\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__25139\,
            I => \N__25136\
        );

    \I__3626\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25133\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__25133\,
            I => \N__25130\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__25130\,
            I => \current_shift_inst.PI_CTRL.integrator_i_3\
        );

    \I__3623\ : InMux
    port map (
            O => \N__25127\,
            I => \N__25124\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__25124\,
            I => \N__25121\
        );

    \I__3621\ : Odrv4
    port map (
            O => \N__25121\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__3620\ : InMux
    port map (
            O => \N__25118\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\
        );

    \I__3619\ : InMux
    port map (
            O => \N__25115\,
            I => \N__25112\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__25112\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__25109\,
            I => \N__25106\
        );

    \I__3616\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25103\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__25103\,
            I => \current_shift_inst.PI_CTRL.integrator_i_4\
        );

    \I__3614\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25097\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__25097\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__3612\ : InMux
    port map (
            O => \N__25094\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\
        );

    \I__3611\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25088\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__25088\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__25085\,
            I => \N__25082\
        );

    \I__3608\ : InMux
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__3606\ : Span4Mux_h
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__3605\ : Odrv4
    port map (
            O => \N__25073\,
            I => \current_shift_inst.PI_CTRL.integrator_i_5\
        );

    \I__3604\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25067\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__25067\,
            I => \N__25064\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__25064\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__3601\ : InMux
    port map (
            O => \N__25061\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\
        );

    \I__3600\ : InMux
    port map (
            O => \N__25058\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\
        );

    \I__3599\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__25052\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__25049\,
            I => \N__25046\
        );

    \I__3596\ : InMux
    port map (
            O => \N__25046\,
            I => \N__25043\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__25043\,
            I => \N__25040\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__25040\,
            I => \current_shift_inst.PI_CTRL.integrator_i_7\
        );

    \I__3593\ : InMux
    port map (
            O => \N__25037\,
            I => \N__25034\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__25034\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3591\ : InMux
    port map (
            O => \N__25031\,
            I => \bfn_10_11_0_\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__25028\,
            I => \N__25025\
        );

    \I__3589\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25021\
        );

    \I__3588\ : InMux
    port map (
            O => \N__25024\,
            I => \N__25018\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__25021\,
            I => \N__25013\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__25018\,
            I => \N__25010\
        );

    \I__3585\ : InMux
    port map (
            O => \N__25017\,
            I => \N__25006\
        );

    \I__3584\ : InMux
    port map (
            O => \N__25016\,
            I => \N__25003\
        );

    \I__3583\ : Span4Mux_h
    port map (
            O => \N__25013\,
            I => \N__25000\
        );

    \I__3582\ : Span4Mux_v
    port map (
            O => \N__25010\,
            I => \N__24997\
        );

    \I__3581\ : InMux
    port map (
            O => \N__25009\,
            I => \N__24994\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__24989\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__25003\,
            I => \N__24989\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__25000\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__24997\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__24994\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__24989\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__24980\,
            I => \N__24977\
        );

    \I__3573\ : InMux
    port map (
            O => \N__24977\,
            I => \N__24973\
        );

    \I__3572\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24970\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__24973\,
            I => \N__24966\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__24970\,
            I => \N__24961\
        );

    \I__3569\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24958\
        );

    \I__3568\ : Span4Mux_h
    port map (
            O => \N__24966\,
            I => \N__24955\
        );

    \I__3567\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24952\
        );

    \I__3566\ : InMux
    port map (
            O => \N__24964\,
            I => \N__24949\
        );

    \I__3565\ : Span4Mux_v
    port map (
            O => \N__24961\,
            I => \N__24944\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__24958\,
            I => \N__24944\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__24955\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__24952\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__24949\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__24944\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3559\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24930\
        );

    \I__3558\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24927\
        );

    \I__3557\ : CascadeMux
    port map (
            O => \N__24933\,
            I => \N__24922\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__24930\,
            I => \N__24919\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__24927\,
            I => \N__24916\
        );

    \I__3554\ : InMux
    port map (
            O => \N__24926\,
            I => \N__24911\
        );

    \I__3553\ : InMux
    port map (
            O => \N__24925\,
            I => \N__24911\
        );

    \I__3552\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24908\
        );

    \I__3551\ : Span4Mux_h
    port map (
            O => \N__24919\,
            I => \N__24905\
        );

    \I__3550\ : Span4Mux_h
    port map (
            O => \N__24916\,
            I => \N__24900\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__24911\,
            I => \N__24900\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__24908\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__24905\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__24900\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__24893\,
            I => \N__24890\
        );

    \I__3544\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24887\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__24887\,
            I => \N__24881\
        );

    \I__3542\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24877\
        );

    \I__3541\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24874\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__24884\,
            I => \N__24871\
        );

    \I__3539\ : Span4Mux_v
    port map (
            O => \N__24881\,
            I => \N__24868\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24865\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__24877\,
            I => \N__24860\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__24874\,
            I => \N__24860\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24857\
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__24868\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__24865\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__24860\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__24857\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__24848\,
            I => \N__24845\
        );

    \I__3529\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24841\
        );

    \I__3528\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24838\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__24841\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_16\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__24838\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_16\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24828\
        );

    \I__3524\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24825\
        );

    \I__3523\ : InMux
    port map (
            O => \N__24831\,
            I => \N__24822\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__24828\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__24825\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__24822\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__3519\ : InMux
    port map (
            O => \N__24815\,
            I => \N__24810\
        );

    \I__3518\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24807\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24804\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__24810\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__24807\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__24804\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__24797\,
            I => \N__24794\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24791\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24791\,
            I => \N__24788\
        );

    \I__3510\ : Span4Mux_v
    port map (
            O => \N__24788\,
            I => \N__24785\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__24785\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__3508\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24779\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24775\
        );

    \I__3506\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24772\
        );

    \I__3505\ : Span4Mux_v
    port map (
            O => \N__24775\,
            I => \N__24768\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__24772\,
            I => \N__24765\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__24771\,
            I => \N__24762\
        );

    \I__3502\ : Span4Mux_h
    port map (
            O => \N__24768\,
            I => \N__24756\
        );

    \I__3501\ : Span4Mux_v
    port map (
            O => \N__24765\,
            I => \N__24756\
        );

    \I__3500\ : InMux
    port map (
            O => \N__24762\,
            I => \N__24751\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24761\,
            I => \N__24751\
        );

    \I__3498\ : Odrv4
    port map (
            O => \N__24756\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24751\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24741\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24738\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__24744\,
            I => \N__24735\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__24741\,
            I => \N__24732\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__24738\,
            I => \N__24729\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24735\,
            I => \N__24724\
        );

    \I__3490\ : Span12Mux_v
    port map (
            O => \N__24732\,
            I => \N__24721\
        );

    \I__3489\ : Span4Mux_v
    port map (
            O => \N__24729\,
            I => \N__24718\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24715\
        );

    \I__3487\ : InMux
    port map (
            O => \N__24727\,
            I => \N__24712\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__24724\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3485\ : Odrv12
    port map (
            O => \N__24721\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3484\ : Odrv4
    port map (
            O => \N__24718\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__24715\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__24712\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__24701\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9_cascade_\
        );

    \I__3480\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24695\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__24695\,
            I => \N__24692\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__24692\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\
        );

    \I__3477\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24683\
        );

    \I__3476\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24683\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__24683\,
            I => \delay_measurement_inst.elapsed_time_hc_28\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24677\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__24677\,
            I => \delay_measurement_inst.N_52\
        );

    \I__3472\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24671\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__3470\ : Glb2LocalMux
    port map (
            O => \N__24668\,
            I => \N__24665\
        );

    \I__3469\ : GlobalMux
    port map (
            O => \N__24665\,
            I => clk_12mhz
        );

    \I__3468\ : IoInMux
    port map (
            O => \N__24662\,
            I => \N__24659\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__24659\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__3466\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24653\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__24653\,
            I => \N__24650\
        );

    \I__3464\ : Span4Mux_h
    port map (
            O => \N__24650\,
            I => \N__24647\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__24647\,
            I => il_min_comp1_c
        );

    \I__3462\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24641\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__3460\ : Span4Mux_h
    port map (
            O => \N__24638\,
            I => \N__24635\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__24635\,
            I => \il_max_comp1_D1\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24629\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__24629\,
            I => \il_min_comp1_D1\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24626\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__3455\ : InMux
    port map (
            O => \N__24623\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__3454\ : InMux
    port map (
            O => \N__24620\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24617\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__3452\ : InMux
    port map (
            O => \N__24614\,
            I => \bfn_9_22_0_\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24611\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__3450\ : InMux
    port map (
            O => \N__24608\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24605\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__3448\ : InMux
    port map (
            O => \N__24602\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__3447\ : CEMux
    port map (
            O => \N__24599\,
            I => \N__24584\
        );

    \I__3446\ : CEMux
    port map (
            O => \N__24598\,
            I => \N__24584\
        );

    \I__3445\ : CEMux
    port map (
            O => \N__24597\,
            I => \N__24584\
        );

    \I__3444\ : CEMux
    port map (
            O => \N__24596\,
            I => \N__24584\
        );

    \I__3443\ : CEMux
    port map (
            O => \N__24595\,
            I => \N__24584\
        );

    \I__3442\ : GlobalMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__3441\ : gio2CtrlBuf
    port map (
            O => \N__24581\,
            I => \delay_measurement_inst.delay_hc_timer.N_302_i_g\
        );

    \I__3440\ : InMux
    port map (
            O => \N__24578\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__3439\ : InMux
    port map (
            O => \N__24575\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__24572\,
            I => \N__24567\
        );

    \I__3437\ : InMux
    port map (
            O => \N__24571\,
            I => \N__24564\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24570\,
            I => \N__24559\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24567\,
            I => \N__24559\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__24564\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__24559\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__3432\ : InMux
    port map (
            O => \N__24554\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24547\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24550\,
            I => \N__24543\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__24547\,
            I => \N__24540\
        );

    \I__3428\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24537\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__24543\,
            I => \N__24534\
        );

    \I__3426\ : Odrv4
    port map (
            O => \N__24540\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__24537\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__3424\ : Odrv4
    port map (
            O => \N__24534\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24527\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__3422\ : InMux
    port map (
            O => \N__24524\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__24521\,
            I => \N__24517\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24520\,
            I => \N__24513\
        );

    \I__3419\ : InMux
    port map (
            O => \N__24517\,
            I => \N__24510\
        );

    \I__3418\ : InMux
    port map (
            O => \N__24516\,
            I => \N__24507\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__24513\,
            I => \N__24502\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__24510\,
            I => \N__24502\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__24507\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__24502\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__3413\ : InMux
    port map (
            O => \N__24497\,
            I => \bfn_9_21_0_\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24494\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__3411\ : InMux
    port map (
            O => \N__24491\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__3410\ : InMux
    port map (
            O => \N__24488\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24481\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24478\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__24481\,
            I => \N__24473\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24473\
        );

    \I__3405\ : Span4Mux_v
    port map (
            O => \N__24473\,
            I => \N__24468\
        );

    \I__3404\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24463\
        );

    \I__3403\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24463\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__24468\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__24463\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__3400\ : InMux
    port map (
            O => \N__24458\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__3399\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24452\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__24452\,
            I => \N__24446\
        );

    \I__3397\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24443\
        );

    \I__3396\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24438\
        );

    \I__3395\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24438\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__24446\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__24443\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__24438\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__3391\ : InMux
    port map (
            O => \N__24431\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__3390\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24424\
        );

    \I__3389\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24421\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__24424\,
            I => \N__24416\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__24421\,
            I => \N__24416\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__24416\,
            I => \N__24411\
        );

    \I__3385\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24408\
        );

    \I__3384\ : InMux
    port map (
            O => \N__24414\,
            I => \N__24405\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__24411\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__24408\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__24405\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24398\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__3379\ : InMux
    port map (
            O => \N__24395\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__3378\ : InMux
    port map (
            O => \N__24392\,
            I => \N__24386\
        );

    \I__3377\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24386\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__24386\,
            I => \N__24382\
        );

    \I__3375\ : InMux
    port map (
            O => \N__24385\,
            I => \N__24379\
        );

    \I__3374\ : Span4Mux_h
    port map (
            O => \N__24382\,
            I => \N__24376\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__24379\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__24376\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__3371\ : InMux
    port map (
            O => \N__24371\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__3370\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24365\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__24365\,
            I => \N__24362\
        );

    \I__3368\ : Span4Mux_h
    port map (
            O => \N__24362\,
            I => \N__24357\
        );

    \I__3367\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24354\
        );

    \I__3366\ : InMux
    port map (
            O => \N__24360\,
            I => \N__24351\
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__24357\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__24354\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__24351\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__3362\ : InMux
    port map (
            O => \N__24344\,
            I => \bfn_9_20_0_\
        );

    \I__3361\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24338\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__24338\,
            I => \N__24333\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__24337\,
            I => \N__24330\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__24336\,
            I => \N__24327\
        );

    \I__3357\ : Span4Mux_v
    port map (
            O => \N__24333\,
            I => \N__24324\
        );

    \I__3356\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24321\
        );

    \I__3355\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24318\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__24324\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__24321\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__24318\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__3351\ : InMux
    port map (
            O => \N__24311\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__3350\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24305\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24300\
        );

    \I__3348\ : InMux
    port map (
            O => \N__24304\,
            I => \N__24295\
        );

    \I__3347\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24295\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__24300\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__24295\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__3344\ : InMux
    port map (
            O => \N__24290\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__3343\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24281\
        );

    \I__3342\ : InMux
    port map (
            O => \N__24286\,
            I => \N__24276\
        );

    \I__3341\ : InMux
    port map (
            O => \N__24285\,
            I => \N__24276\
        );

    \I__3340\ : InMux
    port map (
            O => \N__24284\,
            I => \N__24273\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__24281\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__24276\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__24273\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__24266\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt30_cascade_\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__24263\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1_cascade_\
        );

    \I__3334\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24257\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__24257\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt14_0\
        );

    \I__3332\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24251\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__24251\,
            I => \delay_measurement_inst.N_41\
        );

    \I__3330\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24245\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__24245\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\
        );

    \I__3328\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24235\
        );

    \I__3327\ : InMux
    port map (
            O => \N__24241\,
            I => \N__24235\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24232\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__24235\,
            I => \N__24229\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24224\
        );

    \I__3323\ : Span4Mux_h
    port map (
            O => \N__24229\,
            I => \N__24224\
        );

    \I__3322\ : Odrv4
    port map (
            O => \N__24224\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__3321\ : InMux
    port map (
            O => \N__24221\,
            I => \N__24216\
        );

    \I__3320\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24213\
        );

    \I__3319\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24210\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__24216\,
            I => \N__24207\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__24213\,
            I => \N__24204\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__24210\,
            I => \N__24197\
        );

    \I__3315\ : Span4Mux_v
    port map (
            O => \N__24207\,
            I => \N__24197\
        );

    \I__3314\ : Span4Mux_h
    port map (
            O => \N__24204\,
            I => \N__24197\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__24197\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__3312\ : InMux
    port map (
            O => \N__24194\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__3311\ : InMux
    port map (
            O => \N__24191\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__3310\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24184\
        );

    \I__3309\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24181\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__24184\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__24181\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3306\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24173\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__24173\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__3304\ : InMux
    port map (
            O => \N__24170\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__3303\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24163\
        );

    \I__3302\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24160\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__24163\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__24160\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3299\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24152\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__24152\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__3297\ : InMux
    port map (
            O => \N__24149\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__3296\ : InMux
    port map (
            O => \N__24146\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__3295\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24139\
        );

    \I__3294\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24136\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__24139\,
            I => \N__24133\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__24136\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3291\ : Odrv4
    port map (
            O => \N__24133\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24128\,
            I => \N__24125\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24125\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__3288\ : InMux
    port map (
            O => \N__24122\,
            I => \bfn_9_16_0_\
        );

    \I__3287\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24115\
        );

    \I__3286\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24112\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N__24109\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__24112\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__24109\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3282\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24101\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__24101\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__3280\ : InMux
    port map (
            O => \N__24098\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__3279\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24091\
        );

    \I__3278\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24088\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__24091\,
            I => \N__24085\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__24088\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__24085\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3274\ : InMux
    port map (
            O => \N__24080\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__3273\ : InMux
    port map (
            O => \N__24077\,
            I => \N__24074\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__24074\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__24071\,
            I => \N__24068\
        );

    \I__3270\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24065\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__24065\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__3268\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24058\
        );

    \I__3267\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24055\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__24058\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__24055\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3264\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24047\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__24047\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__3262\ : InMux
    port map (
            O => \N__24044\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__3261\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24037\
        );

    \I__3260\ : InMux
    port map (
            O => \N__24040\,
            I => \N__24034\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__24037\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__24034\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3257\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24026\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__24026\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__3255\ : InMux
    port map (
            O => \N__24023\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__3254\ : InMux
    port map (
            O => \N__24020\,
            I => \N__24016\
        );

    \I__3253\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24013\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24016\,
            I => \N__24010\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__24013\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__24010\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3249\ : InMux
    port map (
            O => \N__24005\,
            I => \N__24002\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__24002\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__3247\ : InMux
    port map (
            O => \N__23999\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__3246\ : InMux
    port map (
            O => \N__23996\,
            I => \N__23992\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23995\,
            I => \N__23989\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__23992\,
            I => \N__23986\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__23989\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__23986\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3241\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__23978\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__3239\ : InMux
    port map (
            O => \N__23975\,
            I => \bfn_9_15_0_\
        );

    \I__3238\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23968\
        );

    \I__3237\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23965\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__23968\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__23965\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3234\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23957\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__23957\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__3232\ : InMux
    port map (
            O => \N__23954\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__3231\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23947\
        );

    \I__3230\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23944\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__23947\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__23944\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3227\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23936\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__23936\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__3225\ : InMux
    port map (
            O => \N__23933\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__3224\ : InMux
    port map (
            O => \N__23930\,
            I => \N__23926\
        );

    \I__3223\ : InMux
    port map (
            O => \N__23929\,
            I => \N__23923\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__23926\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__23923\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3220\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23915\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__23915\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__3218\ : InMux
    port map (
            O => \N__23912\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__3217\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23905\
        );

    \I__3216\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23902\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__23905\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__23902\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3213\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23894\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__23894\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__3211\ : InMux
    port map (
            O => \N__23891\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__3210\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__23885\,
            I => \N__23882\
        );

    \I__3208\ : Span4Mux_h
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__23879\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__23876\,
            I => \N__23873\
        );

    \I__3205\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23869\
        );

    \I__3204\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23865\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__23869\,
            I => \N__23862\
        );

    \I__3202\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23859\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__23865\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__23862\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__23859\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3198\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23848\
        );

    \I__3197\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23845\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__23848\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__23845\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23840\,
            I => \N__23837\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__23837\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__3192\ : InMux
    port map (
            O => \N__23834\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__3191\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23827\
        );

    \I__3190\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23824\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__23827\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__23824\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23816\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__23816\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__3185\ : InMux
    port map (
            O => \N__23813\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__23810\,
            I => \N__23807\
        );

    \I__3183\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23803\
        );

    \I__3182\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23800\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__23803\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__23800\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3179\ : InMux
    port map (
            O => \N__23795\,
            I => \N__23792\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__23792\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__3177\ : InMux
    port map (
            O => \N__23789\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__3176\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23782\
        );

    \I__3175\ : InMux
    port map (
            O => \N__23785\,
            I => \N__23779\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__23782\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__23779\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3172\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23771\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__23771\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__3170\ : InMux
    port map (
            O => \N__23768\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__23765\,
            I => \N__23762\
        );

    \I__3168\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23759\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23759\,
            I => \N__23756\
        );

    \I__3166\ : Span4Mux_v
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__3165\ : Odrv4
    port map (
            O => \N__23753\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__3164\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23747\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__23747\,
            I => \N__23744\
        );

    \I__3162\ : Span4Mux_h
    port map (
            O => \N__23744\,
            I => \N__23739\
        );

    \I__3161\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23736\
        );

    \I__3160\ : InMux
    port map (
            O => \N__23742\,
            I => \N__23733\
        );

    \I__3159\ : Span4Mux_h
    port map (
            O => \N__23739\,
            I => \N__23730\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23727\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__23733\,
            I => \N__23724\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__23730\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__23727\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3154\ : Odrv12
    port map (
            O => \N__23724\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__3152\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23711\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__23711\,
            I => \N__23708\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__23708\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__3149\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23699\
        );

    \I__3148\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23695\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__23703\,
            I => \N__23692\
        );

    \I__3146\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23689\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__23699\,
            I => \N__23686\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23683\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__23695\,
            I => \N__23680\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23677\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__23689\,
            I => \N__23674\
        );

    \I__3140\ : Span4Mux_h
    port map (
            O => \N__23686\,
            I => \N__23667\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__23683\,
            I => \N__23667\
        );

    \I__3138\ : Span4Mux_v
    port map (
            O => \N__23680\,
            I => \N__23667\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__23677\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3136\ : Odrv12
    port map (
            O => \N__23674\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3135\ : Odrv4
    port map (
            O => \N__23667\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23657\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23652\
        );

    \I__3132\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23649\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__23655\,
            I => \N__23645\
        );

    \I__3130\ : Span4Mux_v
    port map (
            O => \N__23652\,
            I => \N__23641\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__23649\,
            I => \N__23638\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23635\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23630\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23644\,
            I => \N__23630\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__23641\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__23638\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__23635\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__23630\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__3118\ : Span4Mux_h
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__3117\ : Odrv4
    port map (
            O => \N__23609\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23600\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__23600\,
            I => \N__23597\
        );

    \I__3113\ : Span4Mux_h
    port map (
            O => \N__23597\,
            I => \N__23594\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__23594\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23587\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23584\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__23587\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__23584\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__3107\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__23576\,
            I => \N__23571\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__23575\,
            I => \N__23568\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__23574\,
            I => \N__23565\
        );

    \I__3103\ : Span12Mux_v
    port map (
            O => \N__23571\,
            I => \N__23561\
        );

    \I__3102\ : InMux
    port map (
            O => \N__23568\,
            I => \N__23558\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23555\
        );

    \I__3100\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23552\
        );

    \I__3099\ : Odrv12
    port map (
            O => \N__23561\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23558\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__23555\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__23552\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__3095\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23538\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23535\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23541\,
            I => \N__23532\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__23538\,
            I => \N__23527\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23535\,
            I => \N__23527\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23532\,
            I => \N__23524\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__23527\,
            I => \N__23521\
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__23524\,
            I => \il_min_comp2_D2\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__23521\,
            I => \il_min_comp2_D2\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23511\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__23515\,
            I => \N__23508\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23514\,
            I => \N__23504\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__23511\,
            I => \N__23501\
        );

    \I__3082\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23496\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23496\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__23504\,
            I => \N__23493\
        );

    \I__3079\ : Span12Mux_v
    port map (
            O => \N__23501\,
            I => \N__23488\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__23496\,
            I => \N__23488\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__23493\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3076\ : Odrv12
    port map (
            O => \N__23488\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__23483\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__3074\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23477\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__23477\,
            I => \current_shift_inst.PI_CTRL.N_72\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__23471\,
            I => \N__23468\
        );

    \I__3070\ : Span4Mux_v
    port map (
            O => \N__23468\,
            I => \N__23465\
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__23465\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__23462\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\
        );

    \I__3067\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23456\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__23456\,
            I => \N__23453\
        );

    \I__3065\ : Odrv4
    port map (
            O => \N__23453\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\
        );

    \I__3064\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__23447\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__23444\,
            I => \delay_measurement_inst.N_30_cascade_\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23438\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__23438\,
            I => \delay_measurement_inst.N_37\
        );

    \I__3059\ : IoInMux
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__23432\,
            I => \N__23429\
        );

    \I__3057\ : Span4Mux_s3_v
    port map (
            O => \N__23429\,
            I => \N__23426\
        );

    \I__3056\ : Span4Mux_v
    port map (
            O => \N__23426\,
            I => \N__23423\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__23423\,
            I => \delay_measurement_inst.delay_hc_timer.N_302_i\
        );

    \I__3054\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23417\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__23417\,
            I => \delay_measurement_inst.N_36\
        );

    \I__3052\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23411\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__23411\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__23408\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9_cascade_\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__23405\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_\
        );

    \I__3048\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__23399\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\
        );

    \I__3046\ : CascadeMux
    port map (
            O => \N__23396\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12_cascade_\
        );

    \I__3045\ : InMux
    port map (
            O => \N__23393\,
            I => \N__23390\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__23390\,
            I => \N__23387\
        );

    \I__3043\ : Odrv12
    port map (
            O => \N__23387\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__23384\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_4_cascade_\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__23378\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__23375\,
            I => \delay_measurement_inst.un1_elapsed_time_hc_cascade_\
        );

    \I__3038\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23369\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__23369\,
            I => \delay_measurement_inst.N_31\
        );

    \I__3036\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23363\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__23363\,
            I => \delay_measurement_inst.N_40\
        );

    \I__3034\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23357\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__23357\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__23354\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_\
        );

    \I__3031\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__23348\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__23345\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1_cascade_\
        );

    \I__3028\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__23339\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt14_0\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__23336\,
            I => \N__23333\
        );

    \I__3025\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__23330\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__3022\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23321\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23318\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__23318\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__3018\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__23309\,
            I => \N__23306\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__23306\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__3014\ : InMux
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__23297\,
            I => \N__23294\
        );

    \I__3012\ : Span4Mux_h
    port map (
            O => \N__23294\,
            I => \N__23291\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__23291\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__23288\,
            I => \N__23285\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23282\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__23282\,
            I => \N__23279\
        );

    \I__3007\ : Span4Mux_v
    port map (
            O => \N__23279\,
            I => \N__23276\
        );

    \I__3006\ : Odrv4
    port map (
            O => \N__23276\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__23273\,
            I => \N__23270\
        );

    \I__3004\ : InMux
    port map (
            O => \N__23270\,
            I => \N__23267\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__23267\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__23264\,
            I => \N__23261\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__2999\ : Span4Mux_v
    port map (
            O => \N__23255\,
            I => \N__23252\
        );

    \I__2998\ : Odrv4
    port map (
            O => \N__23252\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__2997\ : IoInMux
    port map (
            O => \N__23249\,
            I => \N__23246\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__2995\ : Span12Mux_s8_v
    port map (
            O => \N__23243\,
            I => \N__23240\
        );

    \I__2994\ : Odrv12
    port map (
            O => \N__23240\,
            I => s4_phy_c
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__23237\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__23234\,
            I => \N__23231\
        );

    \I__2991\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23228\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__23228\,
            I => \N__23225\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__23225\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__23222\,
            I => \N__23219\
        );

    \I__2987\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__23216\,
            I => \N__23213\
        );

    \I__2985\ : Odrv12
    port map (
            O => \N__23213\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__2984\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23207\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__23207\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__2982\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23201\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__23201\,
            I => \N__23198\
        );

    \I__2980\ : Span4Mux_v
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__2979\ : Odrv4
    port map (
            O => \N__23195\,
            I => \current_shift_inst.PI_CTRL.N_71\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__23192\,
            I => \current_shift_inst.PI_CTRL.N_75_cascade_\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__23189\,
            I => \N__23186\
        );

    \I__2976\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23183\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__23183\,
            I => \N__23180\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__23180\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__23177\,
            I => \N__23174\
        );

    \I__2972\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23171\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__23171\,
            I => \N__23168\
        );

    \I__2970\ : Span4Mux_v
    port map (
            O => \N__23168\,
            I => \N__23165\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__23165\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__23162\,
            I => \N__23159\
        );

    \I__2967\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23156\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__23156\,
            I => \N__23153\
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__23153\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__23150\,
            I => \N__23147\
        );

    \I__2963\ : InMux
    port map (
            O => \N__23147\,
            I => \N__23144\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__23144\,
            I => \N__23141\
        );

    \I__2961\ : Odrv4
    port map (
            O => \N__23141\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__2960\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23135\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__23135\,
            I => \N__23132\
        );

    \I__2958\ : Odrv4
    port map (
            O => \N__23132\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__2957\ : InMux
    port map (
            O => \N__23129\,
            I => \N__23126\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__23126\,
            I => \N__23123\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__23123\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__2954\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__23117\,
            I => \N__23114\
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__23114\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__23111\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__23108\,
            I => \current_shift_inst.PI_CTRL.N_74_cascade_\
        );

    \I__2949\ : InMux
    port map (
            O => \N__23105\,
            I => \N__23102\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__23102\,
            I => \N__23099\
        );

    \I__2947\ : Odrv4
    port map (
            O => \N__23099\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__2946\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23093\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__23093\,
            I => \current_shift_inst.PI_CTRL.un1_enablelt3_0\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__23090\,
            I => \N__23087\
        );

    \I__2943\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23084\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__23084\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\
        );

    \I__2941\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23078\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__23078\,
            I => \delay_measurement_inst.N_32\
        );

    \I__2939\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__23072\,
            I => \delay_measurement_inst.N_35\
        );

    \I__2937\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__23066\,
            I => \N__23063\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__23063\,
            I => \delay_measurement_inst.N_43\
        );

    \I__2934\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23057\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__23057\,
            I => \N__23054\
        );

    \I__2932\ : Odrv12
    port map (
            O => \N__23054\,
            I => il_max_comp1_c
        );

    \I__2931\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23048\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__23048\,
            I => \N__23045\
        );

    \I__2929\ : Span4Mux_v
    port map (
            O => \N__23045\,
            I => \N__23042\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__23042\,
            I => \delay_measurement_inst.N_34\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__23039\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_\
        );

    \I__2926\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23033\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__23033\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__2924\ : InMux
    port map (
            O => \N__23030\,
            I => \N__23027\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__23027\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__2922\ : InMux
    port map (
            O => \N__23024\,
            I => \N__23021\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__23021\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__2920\ : InMux
    port map (
            O => \N__23018\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__23015\,
            I => \N__23012\
        );

    \I__2918\ : InMux
    port map (
            O => \N__23012\,
            I => \N__23009\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__23009\,
            I => \N__23006\
        );

    \I__2916\ : Odrv4
    port map (
            O => \N__23006\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__23003\,
            I => \N__23000\
        );

    \I__2914\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22997\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__22997\,
            I => \N__22994\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__22994\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__22991\,
            I => \N__22988\
        );

    \I__2910\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22985\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__22985\,
            I => \N__22982\
        );

    \I__2908\ : Span4Mux_h
    port map (
            O => \N__22982\,
            I => \N__22979\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__22979\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__2905\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22970\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__22970\,
            I => \N__22967\
        );

    \I__2903\ : Odrv12
    port map (
            O => \N__22967\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\
        );

    \I__2902\ : InMux
    port map (
            O => \N__22964\,
            I => \N__22961\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__22961\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__22958\,
            I => \N__22955\
        );

    \I__2899\ : InMux
    port map (
            O => \N__22955\,
            I => \N__22952\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__22952\,
            I => \N__22949\
        );

    \I__2897\ : Span4Mux_h
    port map (
            O => \N__22949\,
            I => \N__22946\
        );

    \I__2896\ : Span4Mux_h
    port map (
            O => \N__22946\,
            I => \N__22943\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__22943\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__2894\ : InMux
    port map (
            O => \N__22940\,
            I => \N__22937\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__22937\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__22934\,
            I => \N__22931\
        );

    \I__2891\ : InMux
    port map (
            O => \N__22931\,
            I => \N__22928\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__22928\,
            I => \N__22925\
        );

    \I__2889\ : Span4Mux_h
    port map (
            O => \N__22925\,
            I => \N__22922\
        );

    \I__2888\ : Span4Mux_h
    port map (
            O => \N__22922\,
            I => \N__22919\
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__22919\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__2886\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__22913\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__2884\ : InMux
    port map (
            O => \N__22910\,
            I => \N__22907\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__22907\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22901\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__22901\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__2880\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22895\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__22895\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__2878\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22889\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__22889\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__2876\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22883\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__22883\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__2874\ : InMux
    port map (
            O => \N__22880\,
            I => \N__22877\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__22877\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__2872\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22871\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__22871\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__2870\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22865\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__22865\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__2868\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__22859\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22853\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__22853\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__2864\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22847\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__22847\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__2862\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22841\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__22841\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22835\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__22835\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__2858\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22826\
        );

    \I__2857\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22826\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__2855\ : Odrv4
    port map (
            O => \N__22823\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2854\ : InMux
    port map (
            O => \N__22820\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__2853\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22811\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22811\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__22811\,
            I => \N__22808\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__22808\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22805\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2848\ : InMux
    port map (
            O => \N__22802\,
            I => \N__22796\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22801\,
            I => \N__22796\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__22796\,
            I => \N__22793\
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__22793\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22790\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2843\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22783\
        );

    \I__2842\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22780\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__22783\,
            I => \N__22775\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22775\
        );

    \I__2839\ : Span4Mux_h
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__22772\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22769\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22763\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__22763\,
            I => \N__22759\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22756\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__22759\,
            I => \N__22751\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__22756\,
            I => \N__22751\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__22751\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22748\,
            I => \bfn_7_14_0_\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22742\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__22742\,
            I => \N__22738\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22735\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__22738\,
            I => \N__22732\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22729\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__22732\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2823\ : Odrv12
    port map (
            O => \N__22729\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2822\ : InMux
    port map (
            O => \N__22724\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2821\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22717\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22714\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__22717\,
            I => \N__22709\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22714\,
            I => \N__22709\
        );

    \I__2817\ : Odrv4
    port map (
            O => \N__22709\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2816\ : InMux
    port map (
            O => \N__22706\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2815\ : InMux
    port map (
            O => \N__22703\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22700\,
            I => \N__22696\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__22699\,
            I => \N__22693\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__22696\,
            I => \N__22686\
        );

    \I__2811\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22683\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__22692\,
            I => \N__22680\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__22691\,
            I => \N__22677\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__22690\,
            I => \N__22674\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__22689\,
            I => \N__22670\
        );

    \I__2806\ : Span4Mux_s2_h
    port map (
            O => \N__22686\,
            I => \N__22662\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22662\
        );

    \I__2804\ : InMux
    port map (
            O => \N__22680\,
            I => \N__22655\
        );

    \I__2803\ : InMux
    port map (
            O => \N__22677\,
            I => \N__22655\
        );

    \I__2802\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22655\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22652\
        );

    \I__2800\ : InMux
    port map (
            O => \N__22670\,
            I => \N__22649\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22669\,
            I => \N__22646\
        );

    \I__2798\ : InMux
    port map (
            O => \N__22668\,
            I => \N__22641\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22641\
        );

    \I__2796\ : Span4Mux_v
    port map (
            O => \N__22662\,
            I => \N__22638\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__22655\,
            I => \N__22633\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__22652\,
            I => \N__22633\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__22649\,
            I => \N__22626\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__22646\,
            I => \N__22626\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__22641\,
            I => \N__22626\
        );

    \I__2790\ : Span4Mux_v
    port map (
            O => \N__22638\,
            I => \N__22623\
        );

    \I__2789\ : Span4Mux_s3_h
    port map (
            O => \N__22633\,
            I => \N__22620\
        );

    \I__2788\ : Span4Mux_h
    port map (
            O => \N__22626\,
            I => \N__22617\
        );

    \I__2787\ : Span4Mux_h
    port map (
            O => \N__22623\,
            I => \N__22614\
        );

    \I__2786\ : Span4Mux_h
    port map (
            O => \N__22620\,
            I => \N__22611\
        );

    \I__2785\ : Span4Mux_h
    port map (
            O => \N__22617\,
            I => \N__22608\
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__22614\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__22611\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__22608\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__22601\,
            I => \N__22598\
        );

    \I__2780\ : InMux
    port map (
            O => \N__22598\,
            I => \N__22594\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__22597\,
            I => \N__22591\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__22594\,
            I => \N__22588\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22591\,
            I => \N__22585\
        );

    \I__2776\ : Span4Mux_v
    port map (
            O => \N__22588\,
            I => \N__22580\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__22585\,
            I => \N__22580\
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__22580\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2773\ : InMux
    port map (
            O => \N__22577\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22568\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22573\,
            I => \N__22568\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__22565\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22562\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22553\
        );

    \I__2766\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22553\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__22550\,
            I => \N__22547\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__22547\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2762\ : InMux
    port map (
            O => \N__22544\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22534\
        );

    \I__2759\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22531\
        );

    \I__2758\ : Span4Mux_v
    port map (
            O => \N__22534\,
            I => \N__22526\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__22531\,
            I => \N__22526\
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__22526\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2755\ : InMux
    port map (
            O => \N__22523\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2754\ : InMux
    port map (
            O => \N__22520\,
            I => \N__22516\
        );

    \I__2753\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22513\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__22516\,
            I => \N__22510\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__22513\,
            I => \N__22507\
        );

    \I__2750\ : Span4Mux_h
    port map (
            O => \N__22510\,
            I => \N__22502\
        );

    \I__2749\ : Span4Mux_v
    port map (
            O => \N__22507\,
            I => \N__22502\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__22502\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2747\ : InMux
    port map (
            O => \N__22499\,
            I => \bfn_7_13_0_\
        );

    \I__2746\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22490\
        );

    \I__2745\ : InMux
    port map (
            O => \N__22495\,
            I => \N__22490\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__22490\,
            I => \N__22487\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__22487\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22484\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__22481\,
            I => \N__22478\
        );

    \I__2740\ : InMux
    port map (
            O => \N__22478\,
            I => \N__22472\
        );

    \I__2739\ : InMux
    port map (
            O => \N__22477\,
            I => \N__22472\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__2737\ : Span4Mux_h
    port map (
            O => \N__22469\,
            I => \N__22466\
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__22466\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2735\ : InMux
    port map (
            O => \N__22463\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__22460\,
            I => \N__22456\
        );

    \I__2733\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22453\
        );

    \I__2732\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22450\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__22453\,
            I => \N__22445\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__22450\,
            I => \N__22445\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__22445\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2728\ : InMux
    port map (
            O => \N__22442\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__2726\ : InMux
    port map (
            O => \N__22436\,
            I => \N__22433\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__22433\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__2724\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22425\
        );

    \I__2723\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22420\
        );

    \I__2722\ : InMux
    port map (
            O => \N__22428\,
            I => \N__22420\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__22425\,
            I => \N__22415\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__22420\,
            I => \N__22415\
        );

    \I__2719\ : Odrv12
    port map (
            O => \N__22415\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2718\ : InMux
    port map (
            O => \N__22412\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__22409\,
            I => \N__22406\
        );

    \I__2716\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__22403\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2714\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__22394\,
            I => \N__22389\
        );

    \I__2711\ : InMux
    port map (
            O => \N__22393\,
            I => \N__22384\
        );

    \I__2710\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22384\
        );

    \I__2709\ : Sp12to4
    port map (
            O => \N__22389\,
            I => \N__22379\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__22384\,
            I => \N__22379\
        );

    \I__2707\ : Odrv12
    port map (
            O => \N__22379\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2706\ : InMux
    port map (
            O => \N__22376\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__2704\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__22367\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2702\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22360\
        );

    \I__2701\ : InMux
    port map (
            O => \N__22363\,
            I => \N__22357\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__22360\,
            I => \N__22354\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22351\
        );

    \I__2698\ : Span4Mux_h
    port map (
            O => \N__22354\,
            I => \N__22348\
        );

    \I__2697\ : Span4Mux_h
    port map (
            O => \N__22351\,
            I => \N__22345\
        );

    \I__2696\ : Odrv4
    port map (
            O => \N__22348\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__22345\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2694\ : InMux
    port map (
            O => \N__22340\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__22337\,
            I => \N__22333\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__22336\,
            I => \N__22330\
        );

    \I__2691\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22327\
        );

    \I__2690\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22324\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__22327\,
            I => \N__22321\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22318\
        );

    \I__2687\ : Span4Mux_h
    port map (
            O => \N__22321\,
            I => \N__22315\
        );

    \I__2686\ : Span4Mux_h
    port map (
            O => \N__22318\,
            I => \N__22312\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__22315\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__22312\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2683\ : InMux
    port map (
            O => \N__22307\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2682\ : InMux
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__22298\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2679\ : InMux
    port map (
            O => \N__22295\,
            I => \N__22291\
        );

    \I__2678\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22288\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__22291\,
            I => \N__22285\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__22288\,
            I => \N__22282\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__22285\,
            I => \N__22279\
        );

    \I__2674\ : Odrv12
    port map (
            O => \N__22282\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__22279\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2672\ : InMux
    port map (
            O => \N__22274\,
            I => \bfn_7_12_0_\
        );

    \I__2671\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22265\
        );

    \I__2670\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22265\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__22265\,
            I => \N__22262\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__22262\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2667\ : InMux
    port map (
            O => \N__22259\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2666\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22250\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22250\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__22247\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2662\ : InMux
    port map (
            O => \N__22244\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2661\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22235\
        );

    \I__2660\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22235\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__22235\,
            I => \N__22232\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__22232\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2657\ : InMux
    port map (
            O => \N__22229\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__22226\,
            I => \N__22223\
        );

    \I__2655\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__22220\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__22217\,
            I => \N__22213\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__22216\,
            I => \N__22210\
        );

    \I__2651\ : InMux
    port map (
            O => \N__22213\,
            I => \N__22205\
        );

    \I__2650\ : InMux
    port map (
            O => \N__22210\,
            I => \N__22198\
        );

    \I__2649\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22198\
        );

    \I__2648\ : InMux
    port map (
            O => \N__22208\,
            I => \N__22198\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__22205\,
            I => \N__22195\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__22198\,
            I => \N__22192\
        );

    \I__2645\ : Span4Mux_v
    port map (
            O => \N__22195\,
            I => \N__22187\
        );

    \I__2644\ : Span4Mux_v
    port map (
            O => \N__22192\,
            I => \N__22187\
        );

    \I__2643\ : Span4Mux_h
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__22184\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2641\ : InMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__22178\,
            I => \N__22173\
        );

    \I__2639\ : InMux
    port map (
            O => \N__22177\,
            I => \N__22168\
        );

    \I__2638\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22168\
        );

    \I__2637\ : Span12Mux_s2_h
    port map (
            O => \N__22173\,
            I => \N__22163\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__22168\,
            I => \N__22163\
        );

    \I__2635\ : Odrv12
    port map (
            O => \N__22163\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2634\ : InMux
    port map (
            O => \N__22160\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2633\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22152\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22147\
        );

    \I__2631\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22147\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__22152\,
            I => \N__22142\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__22147\,
            I => \N__22142\
        );

    \I__2628\ : Odrv12
    port map (
            O => \N__22142\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2627\ : InMux
    port map (
            O => \N__22139\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2626\ : InMux
    port map (
            O => \N__22136\,
            I => \N__22133\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__22133\,
            I => \N__22128\
        );

    \I__2624\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22123\
        );

    \I__2623\ : InMux
    port map (
            O => \N__22131\,
            I => \N__22123\
        );

    \I__2622\ : Span12Mux_s7_h
    port map (
            O => \N__22128\,
            I => \N__22120\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__22123\,
            I => \N__22117\
        );

    \I__2620\ : Odrv12
    port map (
            O => \N__22120\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2619\ : Odrv12
    port map (
            O => \N__22117\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2618\ : InMux
    port map (
            O => \N__22112\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2617\ : InMux
    port map (
            O => \N__22109\,
            I => \N__22106\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__22106\,
            I => \N__22103\
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__22103\,
            I => il_min_comp2_c
        );

    \I__2614\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__22094\,
            I => \il_min_comp2_D1\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__22091\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__22088\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__22085\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__22082\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\
        );

    \I__2607\ : InMux
    port map (
            O => \N__22079\,
            I => \N__22076\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__22076\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2605\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__22070\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2603\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__22064\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2601\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__22055\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__22052\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_\
        );

    \I__2597\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__22046\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2595\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22040\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__22040\,
            I => \N__22031\
        );

    \I__2593\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22024\
        );

    \I__2592\ : InMux
    port map (
            O => \N__22038\,
            I => \N__22024\
        );

    \I__2591\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22024\
        );

    \I__2590\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22019\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22019\
        );

    \I__2588\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22016\
        );

    \I__2587\ : Span4Mux_v
    port map (
            O => \N__22031\,
            I => \N__22011\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__22024\,
            I => \N__22011\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__22006\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__22016\,
            I => \N__22006\
        );

    \I__2583\ : Span4Mux_h
    port map (
            O => \N__22011\,
            I => \N__22003\
        );

    \I__2582\ : Span4Mux_h
    port map (
            O => \N__22006\,
            I => \N__22000\
        );

    \I__2581\ : Odrv4
    port map (
            O => \N__22003\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__22000\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__21992\,
            I => \N__21989\
        );

    \I__2577\ : Span4Mux_v
    port map (
            O => \N__21989\,
            I => \N__21986\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__21986\,
            I => \il_max_comp2_D1\
        );

    \I__2575\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__2573\ : Odrv12
    port map (
            O => \N__21977\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__2570\ : Span4Mux_s3_h
    port map (
            O => \N__21968\,
            I => \N__21965\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__21965\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2568\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21959\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__21959\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__2565\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__21950\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__21947\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__2562\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__21941\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__2559\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21932\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__2556\ : Odrv4
    port map (
            O => \N__21926\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__2555\ : InMux
    port map (
            O => \N__21923\,
            I => \N__21918\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21915\
        );

    \I__2553\ : InMux
    port map (
            O => \N__21921\,
            I => \N__21912\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__21918\,
            I => \N__21909\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__21915\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__21912\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__21909\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2548\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__21899\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2546\ : InMux
    port map (
            O => \N__21896\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2545\ : IoInMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__2543\ : Span12Mux_s9_v
    port map (
            O => \N__21887\,
            I => \N__21884\
        );

    \I__2542\ : Span12Mux_h
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__2541\ : Odrv12
    port map (
            O => \N__21881\,
            I => pwm_output_c
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__21878\,
            I => \N__21874\
        );

    \I__2539\ : InMux
    port map (
            O => \N__21877\,
            I => \N__21864\
        );

    \I__2538\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21859\
        );

    \I__2537\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21859\
        );

    \I__2536\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21854\
        );

    \I__2535\ : InMux
    port map (
            O => \N__21871\,
            I => \N__21854\
        );

    \I__2534\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21847\
        );

    \I__2533\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21847\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21847\
        );

    \I__2531\ : InMux
    port map (
            O => \N__21867\,
            I => \N__21844\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__21864\,
            I => \N__21841\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__21859\,
            I => \N__21836\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__21854\,
            I => \N__21836\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21831\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__21844\,
            I => \N__21831\
        );

    \I__2525\ : Span4Mux_h
    port map (
            O => \N__21841\,
            I => \N__21828\
        );

    \I__2524\ : Span4Mux_h
    port map (
            O => \N__21836\,
            I => \N__21825\
        );

    \I__2523\ : Span4Mux_h
    port map (
            O => \N__21831\,
            I => \N__21822\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__21828\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__21825\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__21822\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__21815\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__21809\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2516\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__21803\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__2513\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__2511\ : Odrv12
    port map (
            O => \N__21791\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__2510\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__21782\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__21767\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__2502\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__2500\ : Odrv12
    port map (
            O => \N__21758\,
            I => il_max_comp2_c
        );

    \I__2499\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__21752\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21749\,
            I => \N__21744\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21748\,
            I => \N__21741\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21738\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__21744\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__21741\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__21738\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__21728\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21719\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__2486\ : Odrv4
    port map (
            O => \N__21716\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__2485\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21708\
        );

    \I__2484\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21705\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21702\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__21708\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__21705\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__21702\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2479\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21692\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__21692\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__21689\,
            I => \N__21686\
        );

    \I__2476\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21683\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__21683\,
            I => \N__21680\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__21677\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21669\
        );

    \I__2471\ : InMux
    port map (
            O => \N__21673\,
            I => \N__21666\
        );

    \I__2470\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21663\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__21669\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__21666\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__21663\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2466\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__21653\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__21644\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__2461\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21636\
        );

    \I__2460\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21633\
        );

    \I__2459\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21630\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21636\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__21633\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__21630\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2455\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21620\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__21620\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2453\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21612\
        );

    \I__2452\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21609\
        );

    \I__2451\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21606\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__21612\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__21609\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__21606\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__21599\,
            I => \N__21596\
        );

    \I__2446\ : InMux
    port map (
            O => \N__21596\,
            I => \N__21593\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__21593\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__2444\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21587\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__21587\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21581\,
            I => \N__21578\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__21578\,
            I => \N__21575\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__21575\,
            I => \N__21572\
        );

    \I__2438\ : Odrv4
    port map (
            O => \N__21572\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21564\
        );

    \I__2436\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21561\
        );

    \I__2435\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21558\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__21564\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__21561\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__21558\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2431\ : InMux
    port map (
            O => \N__21551\,
            I => \N__21548\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__21548\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__21545\,
            I => \N__21542\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21539\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__21539\,
            I => \N__21536\
        );

    \I__2426\ : Span4Mux_h
    port map (
            O => \N__21536\,
            I => \N__21533\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__21533\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__2424\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21525\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21522\
        );

    \I__2422\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21519\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__21525\,
            I => \N__21516\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__21522\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__21519\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__21516\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2417\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21506\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__21506\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21503\,
            I => \N__21500\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__21500\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__2413\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21494\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__2411\ : Odrv12
    port map (
            O => \N__21491\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21488\,
            I => \N__21485\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__21485\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__2408\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21476\
        );

    \I__2406\ : Span4Mux_v
    port map (
            O => \N__21476\,
            I => \N__21473\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__21473\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21467\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__21467\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21464\,
            I => \N__21461\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__21461\,
            I => \N__21458\
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__21458\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__2399\ : InMux
    port map (
            O => \N__21455\,
            I => \N__21452\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__21452\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__2397\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21446\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__21446\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__2395\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21440\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__2393\ : Odrv12
    port map (
            O => \N__21437\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2392\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21431\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__21431\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__21425\,
            I => \N__21422\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__21422\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__21419\,
            I => \N__21415\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__21418\,
            I => \N__21412\
        );

    \I__2385\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21399\
        );

    \I__2384\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21399\
        );

    \I__2383\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21396\
        );

    \I__2382\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21391\
        );

    \I__2381\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21391\
        );

    \I__2380\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21388\
        );

    \I__2379\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21379\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21379\
        );

    \I__2377\ : InMux
    port map (
            O => \N__21405\,
            I => \N__21379\
        );

    \I__2376\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21379\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__21399\,
            I => \N__21372\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__21396\,
            I => \N__21372\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__21391\,
            I => \N__21372\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__21388\,
            I => \N__21369\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__21379\,
            I => \N__21364\
        );

    \I__2370\ : Span4Mux_v
    port map (
            O => \N__21372\,
            I => \N__21364\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__21369\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2368\ : Odrv4
    port map (
            O => \N__21364\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2367\ : CascadeMux
    port map (
            O => \N__21359\,
            I => \N__21352\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__21358\,
            I => \N__21349\
        );

    \I__2365\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21343\
        );

    \I__2364\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21334\
        );

    \I__2363\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21334\
        );

    \I__2362\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21334\
        );

    \I__2361\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21334\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__21348\,
            I => \N__21331\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__21347\,
            I => \N__21327\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__21346\,
            I => \N__21324\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__21343\,
            I => \N__21318\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__21334\,
            I => \N__21318\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21311\
        );

    \I__2354\ : InMux
    port map (
            O => \N__21330\,
            I => \N__21311\
        );

    \I__2353\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21311\
        );

    \I__2352\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21308\
        );

    \I__2351\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21305\
        );

    \I__2350\ : Span4Mux_v
    port map (
            O => \N__21318\,
            I => \N__21298\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__21311\,
            I => \N__21298\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__21308\,
            I => \N__21298\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21295\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__21298\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__21295\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__21290\,
            I => \N__21283\
        );

    \I__2343\ : InMux
    port map (
            O => \N__21289\,
            I => \N__21274\
        );

    \I__2342\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21274\
        );

    \I__2341\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21274\
        );

    \I__2340\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21274\
        );

    \I__2339\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21270\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__21274\,
            I => \N__21266\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__21273\,
            I => \N__21258\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__21270\,
            I => \N__21255\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__21269\,
            I => \N__21241\
        );

    \I__2334\ : Span4Mux_h
    port map (
            O => \N__21266\,
            I => \N__21238\
        );

    \I__2333\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21233\
        );

    \I__2332\ : InMux
    port map (
            O => \N__21264\,
            I => \N__21233\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21263\,
            I => \N__21226\
        );

    \I__2330\ : InMux
    port map (
            O => \N__21262\,
            I => \N__21226\
        );

    \I__2329\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21226\
        );

    \I__2328\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21223\
        );

    \I__2327\ : Span4Mux_v
    port map (
            O => \N__21255\,
            I => \N__21220\
        );

    \I__2326\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21213\
        );

    \I__2325\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21213\
        );

    \I__2324\ : InMux
    port map (
            O => \N__21252\,
            I => \N__21213\
        );

    \I__2323\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21196\
        );

    \I__2322\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21196\
        );

    \I__2321\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21196\
        );

    \I__2320\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21196\
        );

    \I__2319\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21196\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21196\
        );

    \I__2317\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21196\
        );

    \I__2316\ : InMux
    port map (
            O => \N__21244\,
            I => \N__21196\
        );

    \I__2315\ : InMux
    port map (
            O => \N__21241\,
            I => \N__21193\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__21238\,
            I => \N__21186\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__21233\,
            I => \N__21186\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21186\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__21223\,
            I => \N__21179\
        );

    \I__2310\ : Sp12to4
    port map (
            O => \N__21220\,
            I => \N__21179\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__21213\,
            I => \N__21179\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__21196\,
            I => \N__21167\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__21193\,
            I => \N__21164\
        );

    \I__2306\ : Span4Mux_s2_h
    port map (
            O => \N__21186\,
            I => \N__21161\
        );

    \I__2305\ : Span12Mux_h
    port map (
            O => \N__21179\,
            I => \N__21158\
        );

    \I__2304\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21155\
        );

    \I__2303\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21152\
        );

    \I__2302\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21137\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21175\,
            I => \N__21137\
        );

    \I__2300\ : InMux
    port map (
            O => \N__21174\,
            I => \N__21137\
        );

    \I__2299\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21137\
        );

    \I__2298\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21137\
        );

    \I__2297\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21137\
        );

    \I__2296\ : InMux
    port map (
            O => \N__21170\,
            I => \N__21137\
        );

    \I__2295\ : Span4Mux_s1_h
    port map (
            O => \N__21167\,
            I => \N__21134\
        );

    \I__2294\ : Span4Mux_v
    port map (
            O => \N__21164\,
            I => \N__21129\
        );

    \I__2293\ : Span4Mux_v
    port map (
            O => \N__21161\,
            I => \N__21129\
        );

    \I__2292\ : Odrv12
    port map (
            O => \N__21158\,
            I => \N_19_1\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__21155\,
            I => \N_19_1\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__21152\,
            I => \N_19_1\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__21137\,
            I => \N_19_1\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__21134\,
            I => \N_19_1\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__21129\,
            I => \N_19_1\
        );

    \I__2286\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__21113\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__21110\,
            I => \N__21107\
        );

    \I__2283\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21104\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__2281\ : Span4Mux_h
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__21098\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__2279\ : InMux
    port map (
            O => \N__21095\,
            I => \N__21090\
        );

    \I__2278\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21087\
        );

    \I__2277\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21084\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__21090\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__21087\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__21084\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2273\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21074\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__21074\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2271\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21066\
        );

    \I__2270\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21063\
        );

    \I__2269\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21060\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__21066\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__21063\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__21060\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__21053\,
            I => \N__21050\
        );

    \I__2264\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__2262\ : Span4Mux_s3_h
    port map (
            O => \N__21044\,
            I => \N__21041\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__21041\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2260\ : InMux
    port map (
            O => \N__21038\,
            I => \N__21034\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21030\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__21034\,
            I => \N__21027\
        );

    \I__2257\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21024\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__21030\,
            I => \N__21017\
        );

    \I__2255\ : Span4Mux_h
    port map (
            O => \N__21027\,
            I => \N__21017\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__21024\,
            I => \N__21017\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__21017\,
            I => pwm_duty_input_7
        );

    \I__2252\ : InMux
    port map (
            O => \N__21014\,
            I => \N__21011\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__21011\,
            I => \N__21007\
        );

    \I__2250\ : InMux
    port map (
            O => \N__21010\,
            I => \N__21003\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__21007\,
            I => \N__21000\
        );

    \I__2248\ : InMux
    port map (
            O => \N__21006\,
            I => \N__20997\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__21003\,
            I => pwm_duty_input_5
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__21000\,
            I => pwm_duty_input_5
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__20997\,
            I => pwm_duty_input_5
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__2243\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__20984\,
            I => \N__20981\
        );

    \I__2241\ : Odrv12
    port map (
            O => \N__20981\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\
        );

    \I__2240\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__20975\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__2238\ : InMux
    port map (
            O => \N__20972\,
            I => \N__20969\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__20966\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__2235\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__20960\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__2233\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__20951\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20948\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__2229\ : InMux
    port map (
            O => \N__20945\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__2228\ : InMux
    port map (
            O => \N__20942\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__2227\ : InMux
    port map (
            O => \N__20939\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20936\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__2225\ : InMux
    port map (
            O => \N__20933\,
            I => \bfn_3_10_0_\
        );

    \I__2224\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20916\
        );

    \I__2223\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20916\
        );

    \I__2222\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20916\
        );

    \I__2221\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20916\
        );

    \I__2220\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20909\
        );

    \I__2219\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20906\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20903\
        );

    \I__2217\ : InMux
    port map (
            O => \N__20915\,
            I => \N__20894\
        );

    \I__2216\ : InMux
    port map (
            O => \N__20914\,
            I => \N__20894\
        );

    \I__2215\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20894\
        );

    \I__2214\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20894\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__20909\,
            I => \N__20889\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__20906\,
            I => \N__20889\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__20903\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__20894\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__20889\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2208\ : InMux
    port map (
            O => \N__20882\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__2206\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__20873\,
            I => \N__20869\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20866\
        );

    \I__2203\ : Span4Mux_s2_h
    port map (
            O => \N__20869\,
            I => \N__20863\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20860\
        );

    \I__2201\ : Odrv4
    port map (
            O => \N__20863\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__2200\ : Odrv12
    port map (
            O => \N__20860\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20850\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__20854\,
            I => \N__20847\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20853\,
            I => \N__20844\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20841\
        );

    \I__2195\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20838\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__20844\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__20841\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__20838\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__20831\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__2190\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20825\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__20825\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__20822\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20819\,
            I => \bfn_3_9_0_\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20816\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20813\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__2182\ : Span4Mux_h
    port map (
            O => \N__20804\,
            I => \N__20801\
        );

    \I__2181\ : Span4Mux_v
    port map (
            O => \N__20801\,
            I => \N__20798\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__20798\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20795\,
            I => \bfn_2_17_0_\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20789\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__20789\,
            I => \N__20786\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__20786\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__2172\ : Odrv12
    port map (
            O => \N__20774\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__2171\ : InMux
    port map (
            O => \N__20771\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20764\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20761\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20758\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__20761\,
            I => \N__20755\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__20758\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__2165\ : Odrv12
    port map (
            O => \N__20755\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__2164\ : InMux
    port map (
            O => \N__20750\,
            I => \N__20745\
        );

    \I__2163\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20742\
        );

    \I__2162\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20739\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__20745\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__20742\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__20739\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2158\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20728\
        );

    \I__2157\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20725\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__20728\,
            I => \N__20722\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__20725\,
            I => \N__20719\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__20722\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__2153\ : Odrv12
    port map (
            O => \N__20719\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20709\
        );

    \I__2151\ : InMux
    port map (
            O => \N__20713\,
            I => \N__20706\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20712\,
            I => \N__20703\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__20709\,
            I => \N__20700\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__20706\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__20703\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__20700\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20689\
        );

    \I__2144\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20686\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__20689\,
            I => \N__20683\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__20686\,
            I => \N__20680\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__20683\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__2140\ : Odrv12
    port map (
            O => \N__20680\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__20672\,
            I => \N__20668\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20671\,
            I => \N__20664\
        );

    \I__2136\ : Span4Mux_s2_h
    port map (
            O => \N__20668\,
            I => \N__20661\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20658\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__20664\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__20661\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__20658\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2131\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20647\
        );

    \I__2130\ : InMux
    port map (
            O => \N__20650\,
            I => \N__20644\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20647\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__20644\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2127\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20633\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20633\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__2124\ : Odrv12
    port map (
            O => \N__20630\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2123\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20624\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__20624\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__20621\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\
        );

    \I__2120\ : InMux
    port map (
            O => \N__20618\,
            I => \N__20613\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__20617\,
            I => \N__20608\
        );

    \I__2118\ : InMux
    port map (
            O => \N__20616\,
            I => \N__20605\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__20613\,
            I => \N__20602\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20593\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20590\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20587\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__20605\,
            I => \N__20582\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__20602\,
            I => \N__20582\
        );

    \I__2111\ : InMux
    port map (
            O => \N__20601\,
            I => \N__20579\
        );

    \I__2110\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20568\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20568\
        );

    \I__2108\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20568\
        );

    \I__2107\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20568\
        );

    \I__2106\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20568\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__20593\,
            I => \N__20565\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__20590\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__20587\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__20582\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__20579\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20568\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2099\ : Odrv12
    port map (
            O => \N__20565\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__20546\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20543\,
            I => \N__20540\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20540\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__2093\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20534\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__20534\,
            I => \N__20531\
        );

    \I__2091\ : Odrv4
    port map (
            O => \N__20531\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__2090\ : InMux
    port map (
            O => \N__20528\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20522\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__20522\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20519\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__20516\,
            I => \N__20513\
        );

    \I__2085\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20510\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__20510\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20507\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20501\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__20501\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__2080\ : InMux
    port map (
            O => \N__20498\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__2079\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20492\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__20492\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20489\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20483\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20483\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__2074\ : InMux
    port map (
            O => \N__20480\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__2073\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20474\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__20474\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20471\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__2070\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20465\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__20465\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__2068\ : InMux
    port map (
            O => \N__20462\,
            I => \N__20459\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__20459\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__2066\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20453\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__20453\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__2064\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20447\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__20447\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__2062\ : InMux
    port map (
            O => \N__20444\,
            I => \N__20441\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__20441\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__2060\ : InMux
    port map (
            O => \N__20438\,
            I => \N__20435\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__20435\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__2058\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__20429\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__2056\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__20423\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__2054\ : InMux
    port map (
            O => \N__20420\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__2052\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__20411\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__2050\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__20405\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__2048\ : InMux
    port map (
            O => \N__20402\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__2046\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__20393\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__2044\ : InMux
    port map (
            O => \N__20390\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__2043\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20384\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__20384\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__2041\ : InMux
    port map (
            O => \N__20381\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__2040\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__20375\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__2038\ : InMux
    port map (
            O => \N__20372\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__2037\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20366\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__20366\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__2035\ : InMux
    port map (
            O => \N__20363\,
            I => \bfn_2_14_0_\
        );

    \I__2034\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__20357\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__2032\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__20351\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__2030\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__20345\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__20342\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__2027\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20334\
        );

    \I__2026\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20329\
        );

    \I__2025\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20329\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__20334\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__20329\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__20324\,
            I => \N__20320\
        );

    \I__2021\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20316\
        );

    \I__2020\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20313\
        );

    \I__2019\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20310\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__20316\,
            I => \N__20307\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__20313\,
            I => \N__20302\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__20310\,
            I => \N__20302\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__20307\,
            I => pwm_duty_input_9
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__20302\,
            I => pwm_duty_input_9
        );

    \I__2013\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20292\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20289\
        );

    \I__2011\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20286\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__20292\,
            I => pwm_duty_input_6
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__20289\,
            I => pwm_duty_input_6
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__20286\,
            I => pwm_duty_input_6
        );

    \I__2007\ : InMux
    port map (
            O => \N__20279\,
            I => \N__20276\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__20273\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__20270\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\
        );

    \I__2003\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20262\
        );

    \I__2002\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20259\
        );

    \I__2001\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20256\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__20262\,
            I => pwm_duty_input_8
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__20259\,
            I => pwm_duty_input_8
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__20256\,
            I => pwm_duty_input_8
        );

    \I__1997\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20244\
        );

    \I__1996\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20239\
        );

    \I__1995\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20239\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__20244\,
            I => \N__20236\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__20239\,
            I => \N__20233\
        );

    \I__1992\ : Span4Mux_s1_h
    port map (
            O => \N__20236\,
            I => \N__20230\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__20233\,
            I => pwm_duty_input_3
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__20230\,
            I => pwm_duty_input_3
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__20225\,
            I => \N__20222\
        );

    \I__1988\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__20219\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20210\
        );

    \I__1985\ : InMux
    port map (
            O => \N__20215\,
            I => \N__20210\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__20210\,
            I => \N__20206\
        );

    \I__1983\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20203\
        );

    \I__1982\ : Span4Mux_h
    port map (
            O => \N__20206\,
            I => \N__20198\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__20203\,
            I => \N__20198\
        );

    \I__1980\ : Span4Mux_s1_h
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__20195\,
            I => pwm_duty_input_4
        );

    \I__1978\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20188\
        );

    \I__1977\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20185\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__20188\,
            I => \N__20182\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__20185\,
            I => \N__20179\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__20182\,
            I => \N__20176\
        );

    \I__1973\ : Span4Mux_v
    port map (
            O => \N__20179\,
            I => \N__20173\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__20176\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__20173\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1970\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20165\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__20165\,
            I => \N__20162\
        );

    \I__1968\ : Span4Mux_h
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__20159\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1966\ : InMux
    port map (
            O => \N__20156\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1965\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__20150\,
            I => \N__20147\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__20144\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1961\ : InMux
    port map (
            O => \N__20141\,
            I => \N__20138\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__20138\,
            I => \N__20135\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__20135\,
            I => \N__20131\
        );

    \I__1958\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20128\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__20131\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__20128\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__1955\ : InMux
    port map (
            O => \N__20123\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1954\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__20111\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1950\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20105\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__20105\,
            I => \N__20101\
        );

    \I__1948\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20098\
        );

    \I__1947\ : Span4Mux_s2_h
    port map (
            O => \N__20101\,
            I => \N__20093\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__20098\,
            I => \N__20093\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__20093\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1944\ : InMux
    port map (
            O => \N__20090\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__20087\,
            I => \current_shift_inst.PI_CTRL.N_168_cascade_\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__20084\,
            I => \N__20079\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__20083\,
            I => \N__20076\
        );

    \I__1940\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20066\
        );

    \I__1939\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20066\
        );

    \I__1938\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20066\
        );

    \I__1937\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20066\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__20066\,
            I => \current_shift_inst.PI_CTRL.N_166\
        );

    \I__1935\ : InMux
    port map (
            O => \N__20063\,
            I => \N__20059\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20055\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__20059\,
            I => \N__20052\
        );

    \I__1932\ : InMux
    port map (
            O => \N__20058\,
            I => \N__20049\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__20055\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__20052\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__20049\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__1928\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__20039\,
            I => \N__20035\
        );

    \I__1926\ : InMux
    port map (
            O => \N__20038\,
            I => \N__20032\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__20035\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__20032\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__20027\,
            I => \current_shift_inst.PI_CTRL.N_166_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20015\
        );

    \I__1921\ : InMux
    port map (
            O => \N__20023\,
            I => \N__20015\
        );

    \I__1920\ : InMux
    port map (
            O => \N__20022\,
            I => \N__20015\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__20015\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1918\ : InMux
    port map (
            O => \N__20012\,
            I => \N__20009\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__20009\,
            I => \current_shift_inst.PI_CTRL.N_162\
        );

    \I__1916\ : InMux
    port map (
            O => \N__20006\,
            I => \N__20002\
        );

    \I__1915\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19999\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20002\,
            I => \N__19996\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__19999\,
            I => pwm_duty_input_0
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__19996\,
            I => pwm_duty_input_0
        );

    \I__1911\ : InMux
    port map (
            O => \N__19991\,
            I => \N__19987\
        );

    \I__1910\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19984\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__19987\,
            I => \N__19981\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__19984\,
            I => pwm_duty_input_1
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__19981\,
            I => pwm_duty_input_1
        );

    \I__1906\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19972\
        );

    \I__1905\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19969\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__19972\,
            I => \N__19966\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__19969\,
            I => pwm_duty_input_2
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__19966\,
            I => pwm_duty_input_2
        );

    \I__1901\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19952\
        );

    \I__1900\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19952\
        );

    \I__1899\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19952\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__19952\,
            I => \current_shift_inst.PI_CTRL.N_167\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__19949\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\
        );

    \I__1896\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19942\
        );

    \I__1895\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19939\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__19942\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__19939\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1892\ : InMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__19928\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__1889\ : InMux
    port map (
            O => \N__19925\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__1888\ : InMux
    port map (
            O => \N__19922\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__1887\ : InMux
    port map (
            O => \N__19919\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__19913\,
            I => \N_34_i_i\
        );

    \I__1884\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__19907\,
            I => \rgb_drv_RNOZ0\
        );

    \I__1882\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__19901\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__1880\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__1878\ : Span4Mux_v
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__19889\,
            I => \N__19886\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__19886\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1875\ : InMux
    port map (
            O => \N__19883\,
            I => \N__19880\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__19880\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__1873\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__19874\,
            I => \N__19870\
        );

    \I__1871\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19867\
        );

    \I__1870\ : Span4Mux_s2_h
    port map (
            O => \N__19870\,
            I => \N__19864\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__19867\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__19864\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1867\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__1865\ : Span4Mux_v
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__19850\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__1863\ : InMux
    port map (
            O => \N__19847\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__1862\ : InMux
    port map (
            O => \N__19844\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__1861\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__19832\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__1857\ : InMux
    port map (
            O => \N__19829\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__1856\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19822\
        );

    \I__1855\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19818\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__19822\,
            I => \N__19815\
        );

    \I__1853\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19812\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__19818\,
            I => \N__19807\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__19815\,
            I => \N__19807\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__19812\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__19807\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__1847\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__19793\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__1844\ : InMux
    port map (
            O => \N__19790\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__1843\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19782\
        );

    \I__1842\ : InMux
    port map (
            O => \N__19786\,
            I => \N__19779\
        );

    \I__1841\ : InMux
    port map (
            O => \N__19785\,
            I => \N__19776\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__19782\,
            I => \N__19773\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__19779\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__19776\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__19773\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__1835\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__1833\ : Odrv12
    port map (
            O => \N__19757\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__1832\ : InMux
    port map (
            O => \N__19754\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__1830\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__1828\ : Odrv12
    port map (
            O => \N__19742\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__1827\ : InMux
    port map (
            O => \N__19739\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__19727\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__1822\ : InMux
    port map (
            O => \N__19724\,
            I => \bfn_1_19_0_\
        );

    \I__1821\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__19709\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1816\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__19703\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__1814\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19697\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__1812\ : Span4Mux_v
    port map (
            O => \N__19694\,
            I => \N__19691\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__19691\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19685\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__19685\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__1808\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__1806\ : Span4Mux_h
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__19670\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__19664\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__19649\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1796\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__19643\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__1794\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__19631\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__19625\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__1788\ : InMux
    port map (
            O => \N__19622\,
            I => \N__19619\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__1786\ : Span4Mux_h
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__19610\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__19604\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__1781\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__19592\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1777\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__19586\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__1775\ : InMux
    port map (
            O => \N__19583\,
            I => \N__19580\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__1773\ : Span4Mux_v
    port map (
            O => \N__19577\,
            I => \N__19574\
        );

    \I__1772\ : Span4Mux_v
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__19571\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1770\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__19565\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__19562\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19553\
        );

    \I__1766\ : InMux
    port map (
            O => \N__19558\,
            I => \N__19553\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__19547\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__19544\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\
        );

    \I__1761\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__1758\ : Span4Mux_v
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__19529\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__19523\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__1754\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19517\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__19517\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__1751\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__1749\ : Span4Mux_v
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__19502\,
            I => \N__19499\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__19499\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1746\ : InMux
    port map (
            O => \N__19496\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__1744\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19487\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__19487\,
            I => \N__19484\
        );

    \I__1742\ : Span4Mux_v
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__19478\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1739\ : InMux
    port map (
            O => \N__19475\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1738\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19469\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__19469\,
            I => \N__19466\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__19466\,
            I => \N__19463\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__19460\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1733\ : InMux
    port map (
            O => \N__19457\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__1731\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19448\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__19448\,
            I => \N__19445\
        );

    \I__1729\ : Span4Mux_v
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__1728\ : Span4Mux_v
    port map (
            O => \N__19442\,
            I => \N__19439\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__19439\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1726\ : InMux
    port map (
            O => \N__19436\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1725\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19430\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__1722\ : Span4Mux_v
    port map (
            O => \N__19424\,
            I => \N__19421\
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__19421\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1720\ : InMux
    port map (
            O => \N__19418\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__1718\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19409\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19406\
        );

    \I__1716\ : Span4Mux_v
    port map (
            O => \N__19406\,
            I => \N__19403\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__19400\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1713\ : InMux
    port map (
            O => \N__19397\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1712\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19391\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__19391\,
            I => \N__19388\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__19382\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1707\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19375\
        );

    \I__1706\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19372\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__19375\,
            I => \N__19369\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__19372\,
            I => \N__19366\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__19369\,
            I => \N__19360\
        );

    \I__1702\ : Span4Mux_h
    port map (
            O => \N__19366\,
            I => \N__19357\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__19365\,
            I => \N__19354\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__19364\,
            I => \N__19350\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__19363\,
            I => \N__19346\
        );

    \I__1698\ : Span4Mux_v
    port map (
            O => \N__19360\,
            I => \N__19342\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__19357\,
            I => \N__19339\
        );

    \I__1696\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19326\
        );

    \I__1695\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19326\
        );

    \I__1694\ : InMux
    port map (
            O => \N__19350\,
            I => \N__19326\
        );

    \I__1693\ : InMux
    port map (
            O => \N__19349\,
            I => \N__19326\
        );

    \I__1692\ : InMux
    port map (
            O => \N__19346\,
            I => \N__19326\
        );

    \I__1691\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19326\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__19342\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__19339\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__19326\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1687\ : InMux
    port map (
            O => \N__19319\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1686\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__19310\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1683\ : InMux
    port map (
            O => \N__19307\,
            I => \bfn_1_15_0_\
        );

    \I__1682\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__19301\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__1679\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__1677\ : Span4Mux_v
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__19283\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19280\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1673\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__19274\,
            I => \N__19271\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__19265\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__19262\,
            I => \N__19259\
        );

    \I__1667\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__19256\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1665\ : InMux
    port map (
            O => \N__19253\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__19247\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__19244\,
            I => \N__19241\
        );

    \I__1661\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__19229\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1656\ : InMux
    port map (
            O => \N__19226\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1655\ : InMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__19220\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__1652\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19211\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__19208\,
            I => \N__19205\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__19202\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1647\ : InMux
    port map (
            O => \N__19199\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1646\ : InMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__19193\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__1643\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__1641\ : Span4Mux_v
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__1640\ : Span4Mux_v
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__19175\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1638\ : InMux
    port map (
            O => \N__19172\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1637\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__19166\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__19163\,
            I => \N__19160\
        );

    \I__1634\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__1632\ : Span4Mux_v
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__19148\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1629\ : InMux
    port map (
            O => \N__19145\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1628\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__19139\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__1625\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__1622\ : Span4Mux_v
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__19121\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1620\ : InMux
    port map (
            O => \N__19118\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1619\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19112\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__19109\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__1615\ : InMux
    port map (
            O => \N__19103\,
            I => \N__19100\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__1612\ : Span4Mux_v
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__19091\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1610\ : InMux
    port map (
            O => \N__19088\,
            I => \bfn_1_14_0_\
        );

    \I__1609\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__19073\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__1603\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__19061\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1600\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19054\
        );

    \I__1599\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19051\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__19054\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__19051\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__1595\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__19040\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_10_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            carryinitout => \bfn_10_11_0_\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            carryinitout => \bfn_10_12_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_15_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_2_0_\
        );

    \IN_MUX_bfv_15_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_15_3_0_\
        );

    \IN_MUX_bfv_15_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_15_4_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_16_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_14_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_3_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_3_10_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_16_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_7_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_15_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_15_27_0_\
        );

    \IN_MUX_bfv_15_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_15_28_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_12_11_0_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__23435\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_302_i_g\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__34529\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_181_i_g\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__29075\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_304_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__45908\,
            CLKHFEN => \N__45912\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__45967\,
            RGB2PWM => \N__19916\,
            RGB1 => rgb_g_wire,
            CURREN => \N__46081\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__19910\,
            RGB0PWM => \N__47925\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__19379\,
            in1 => \N__21177\,
            in2 => \_gnd_net_\,
            in3 => \N__19057\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22700\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48482\,
            ce => 'H',
            sr => \N__47816\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__19058\,
            in1 => \N__19378\,
            in2 => \N__19046\,
            in3 => \N__21178\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__22400\,
            in1 => \N__21877\,
            in2 => \N__22699\,
            in3 => \N__22043\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48480\,
            ce => 'H',
            sr => \N__47841\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001100"
        )
    port map (
            in0 => \N__22036\,
            in1 => \N__22136\,
            in2 => \N__22689\,
            in3 => \N__21873\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__47850\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__19946\,
            in1 => \N__20012\,
            in2 => \N__22217\,
            in3 => \N__22035\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__47850\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__20023\,
            in1 => \N__21974\,
            in2 => \N__20083\,
            in3 => \N__19960\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__47850\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__19959\,
            in1 => \N__20075\,
            in2 => \N__21053\,
            in3 => \N__20022\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__47850\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__20024\,
            in1 => \N__21983\,
            in2 => \N__20084\,
            in3 => \N__19961\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__47850\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011011101"
        )
    port map (
            in0 => \N__20082\,
            in1 => \N__20062\,
            in2 => \N__21878\,
            in3 => \N__20042\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__47850\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__22430\,
            in1 => \N__21870\,
            in2 => \N__22692\,
            in3 => \N__22039\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48474\,
            ce => 'H',
            sr => \N__47856\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__22157\,
            in1 => \N__21869\,
            in2 => \N__22691\,
            in3 => \N__22038\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48474\,
            ce => 'H',
            sr => \N__47856\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__22181\,
            in1 => \N__21868\,
            in2 => \N__22690\,
            in3 => \N__22037\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48474\,
            ce => 'H',
            sr => \N__47856\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20296\,
            in1 => \N__21037\,
            in2 => \N__20324\,
            in3 => \N__21010\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20134\,
            in2 => \_gnd_net_\,
            in3 => \N__19821\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19085\,
            in2 => \N__19070\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19304\,
            in2 => \N__19298\,
            in3 => \N__19280\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19277\,
            in2 => \N__19262\,
            in3 => \N__19253\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19250\,
            in2 => \N__19244\,
            in3 => \N__19226\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19223\,
            in2 => \N__19217\,
            in3 => \N__19199\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19196\,
            in2 => \N__19190\,
            in3 => \N__19172\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19169\,
            in2 => \N__19163\,
            in3 => \N__19145\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19142\,
            in2 => \N__19136\,
            in3 => \N__19118\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19115\,
            in2 => \N__19106\,
            in3 => \N__19088\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19520\,
            in2 => \N__19514\,
            in3 => \N__19496\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19345\,
            in2 => \N__19493\,
            in3 => \N__19475\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19472\,
            in2 => \N__19363\,
            in3 => \N__19457\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19349\,
            in2 => \N__19454\,
            in3 => \N__19436\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19433\,
            in2 => \N__19364\,
            in3 => \N__19418\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19353\,
            in2 => \N__19415\,
            in3 => \N__19397\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19394\,
            in2 => \N__19365\,
            in3 => \N__19319\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19316\,
            in2 => \N__20417\,
            in3 => \N__19307\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__19841\,
            in1 => \N__20693\,
            in2 => \N__19562\,
            in3 => \N__20675\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20104\,
            in2 => \_gnd_net_\,
            in3 => \N__19786\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20141\,
            in1 => \N__19825\,
            in2 => \N__19802\,
            in3 => \N__20601\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20768\,
            in1 => \N__20749\,
            in2 => \N__19751\,
            in3 => \N__20598\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19873\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19558\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19559\,
            in1 => \N__19859\,
            in2 => \N__19544\,
            in3 => \N__20596\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20732\,
            in1 => \N__20712\,
            in2 => \N__19736\,
            in3 => \N__20599\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__20855\,
            in1 => \N__19934\,
            in2 => \N__20879\,
            in3 => \N__20600\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__20597\,
            in1 => \N__20108\,
            in2 => \N__19766\,
            in3 => \N__19785\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19526\,
            in2 => \_gnd_net_\,
            in3 => \N__19541\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19706\,
            in2 => \_gnd_net_\,
            in3 => \N__19721\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19688\,
            in2 => \_gnd_net_\,
            in3 => \N__19700\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19667\,
            in2 => \_gnd_net_\,
            in3 => \N__19682\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19646\,
            in2 => \_gnd_net_\,
            in3 => \N__19661\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19628\,
            in2 => \_gnd_net_\,
            in3 => \N__19640\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19607\,
            in2 => \_gnd_net_\,
            in3 => \N__19622\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19589\,
            in2 => \_gnd_net_\,
            in3 => \N__19601\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19568\,
            in2 => \_gnd_net_\,
            in3 => \N__19583\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19883\,
            in2 => \_gnd_net_\,
            in3 => \N__19898\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19877\,
            in2 => \_gnd_net_\,
            in3 => \N__19847\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__20612\,
            in1 => \N__20192\,
            in2 => \_gnd_net_\,
            in3 => \N__19844\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20667\,
            in2 => \_gnd_net_\,
            in3 => \N__19829\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19826\,
            in2 => \_gnd_net_\,
            in3 => \N__19790\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19787\,
            in2 => \_gnd_net_\,
            in3 => \N__19754\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20748\,
            in2 => \_gnd_net_\,
            in3 => \N__19739\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20714\,
            in2 => \_gnd_net_\,
            in3 => \N__19724\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20854\,
            in3 => \N__19925\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20650\,
            in2 => \_gnd_net_\,
            in3 => \N__19922\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19919\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_0_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45541\,
            in2 => \_gnd_net_\,
            in3 => \N__47923\,
            lcout => \N_34_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__47924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45545\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_8_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19904\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48477\,
            ce => 'H',
            sr => \N__47832\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24746\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48477\,
            ce => 'H',
            sr => \N__47832\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__21323\,
            in1 => \N__21408\,
            in2 => \N__21269\,
            in3 => \N__20810\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48477\,
            ce => 'H',
            sr => \N__47832\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__22209\,
            in1 => \N__22667\,
            in2 => \_gnd_net_\,
            in3 => \N__20337\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22208\,
            in2 => \_gnd_net_\,
            in3 => \N__20058\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__22669\,
            in1 => \N__19945\,
            in2 => \N__20087\,
            in3 => \N__22034\,
            lcout => \current_shift_inst.PI_CTRL.N_166\,
            ltout => \current_shift_inst.PI_CTRL.N_166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010100"
        )
    port map (
            in0 => \N__20063\,
            in1 => \N__20038\,
            in2 => \N__20027\,
            in3 => \N__21871\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__21872\,
            in1 => \N__22668\,
            in2 => \N__22216\,
            in3 => \N__20338\,
            lcout => \current_shift_inst.PI_CTRL.N_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20005\,
            in1 => \N__19990\,
            in2 => \_gnd_net_\,
            in3 => \N__19975\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__22673\,
            in1 => \N__20339\,
            in2 => \_gnd_net_\,
            in3 => \N__21867\,
            lcout => \current_shift_inst.PI_CTRL.N_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__22429\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22176\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22132\,
            in1 => \N__22393\,
            in2 => \N__19949\,
            in3 => \N__22156\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22428\,
            in2 => \_gnd_net_\,
            in3 => \N__22155\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22392\,
            in1 => \N__22131\,
            in2 => \N__20342\,
            in3 => \N__22177\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20266\,
            in1 => \N__20323\,
            in2 => \N__20990\,
            in3 => \N__20297\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__20279\,
            in1 => \N__20247\,
            in2 => \N__20270\,
            in3 => \N__20215\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__20267\,
            in1 => \N__20248\,
            in2 => \N__20225\,
            in3 => \N__20216\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20191\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20168\,
            in2 => \_gnd_net_\,
            in3 => \N__20156\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20153\,
            in2 => \_gnd_net_\,
            in3 => \N__20123\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20120\,
            in2 => \_gnd_net_\,
            in3 => \N__20090\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20408\,
            in2 => \_gnd_net_\,
            in3 => \N__20402\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45836\,
            in2 => \N__20399\,
            in3 => \N__20390\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20387\,
            in2 => \N__45889\,
            in3 => \N__20381\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20378\,
            in2 => \N__45856\,
            in3 => \N__20372\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20369\,
            in2 => \_gnd_net_\,
            in3 => \N__20363\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20360\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20354\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20348\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20468\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20462\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20456\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20450\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20444\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20438\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20432\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20426\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20420\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20543\,
            in2 => \N__20617\,
            in3 => \N__20611\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20537\,
            in2 => \_gnd_net_\,
            in3 => \N__20528\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20525\,
            in2 => \_gnd_net_\,
            in3 => \N__20519\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20516\,
            in3 => \N__20507\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20504\,
            in2 => \_gnd_net_\,
            in3 => \N__20498\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20495\,
            in2 => \_gnd_net_\,
            in3 => \N__20489\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20486\,
            in2 => \_gnd_net_\,
            in3 => \N__20480\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20477\,
            in2 => \_gnd_net_\,
            in3 => \N__20471\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20552\,
            in3 => \N__20795\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__20792\,
            in1 => \N__20616\,
            in2 => \N__20783\,
            in3 => \N__20771\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20750\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20767\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20713\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20731\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20671\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20692\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20651\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20638\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20639\,
            in1 => \N__20627\,
            in2 => \N__20621\,
            in3 => \N__20618\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34008\,
            in1 => \N__34284\,
            in2 => \N__33592\,
            in3 => \N__34183\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48405\,
            ce => \N__28847\,
            sr => \N__47882\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34184\,
            in1 => \N__33703\,
            in2 => \N__34336\,
            in3 => \N__34009\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48405\,
            ce => \N__28847\,
            sr => \N__47882\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20872\,
            in2 => \_gnd_net_\,
            in3 => \N__20853\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNITBL3_9_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21923\,
            in1 => \N__21530\,
            in2 => \_gnd_net_\,
            in3 => \N__21640\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIRPD2_0_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21093\,
            in2 => \_gnd_net_\,
            in3 => \N__21069\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_2_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__21673\,
            in1 => \N__21712\,
            in2 => \N__20831\,
            in3 => \N__21748\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_6_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20828\,
            in1 => \N__21568\,
            in2 => \N__20822\,
            in3 => \N__21617\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20927\,
            in1 => \N__21095\,
            in2 => \_gnd_net_\,
            in3 => \N__20819\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__47823\
        );

    \pwm_generator_inst.counter_1_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20912\,
            in1 => \N__21071\,
            in2 => \_gnd_net_\,
            in3 => \N__20816\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__47823\
        );

    \pwm_generator_inst.counter_2_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20928\,
            in1 => \N__21749\,
            in2 => \_gnd_net_\,
            in3 => \N__20813\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__47823\
        );

    \pwm_generator_inst.counter_3_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20913\,
            in1 => \N__21713\,
            in2 => \_gnd_net_\,
            in3 => \N__20948\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__47823\
        );

    \pwm_generator_inst.counter_4_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20929\,
            in1 => \N__21674\,
            in2 => \_gnd_net_\,
            in3 => \N__20945\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__47823\
        );

    \pwm_generator_inst.counter_5_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20914\,
            in1 => \N__21641\,
            in2 => \_gnd_net_\,
            in3 => \N__20942\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__47823\
        );

    \pwm_generator_inst.counter_6_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20930\,
            in1 => \N__21616\,
            in2 => \_gnd_net_\,
            in3 => \N__20939\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__47823\
        );

    \pwm_generator_inst.counter_7_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20915\,
            in1 => \N__21569\,
            in2 => \_gnd_net_\,
            in3 => \N__20936\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__47823\
        );

    \pwm_generator_inst.counter_8_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20926\,
            in1 => \N__21529\,
            in2 => \_gnd_net_\,
            in3 => \N__20933\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_10_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__48469\,
            ce => 'H',
            sr => \N__47833\
        );

    \pwm_generator_inst.counter_9_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20925\,
            in1 => \N__21922\,
            in2 => \_gnd_net_\,
            in3 => \N__20882\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48469\,
            ce => 'H',
            sr => \N__47833\
        );

    \pwm_generator_inst.threshold_6_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21482\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48469\,
            ce => 'H',
            sr => \N__47833\
        );

    \pwm_generator_inst.threshold_5_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21443\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48469\,
            ce => 'H',
            sr => \N__47833\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23750\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48462\,
            ce => 'H',
            sr => \N__47842\
        );

    \pwm_generator_inst.threshold_3_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21497\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48462\,
            ce => 'H',
            sr => \N__47842\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21038\,
            in2 => \_gnd_net_\,
            in3 => \N__21014\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_0_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20957\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48443\,
            ce => 'H',
            sr => \N__47857\
        );

    \pwm_generator_inst.threshold_7_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20972\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48443\,
            ce => 'H',
            sr => \N__47857\
        );

    \pwm_generator_inst.threshold_9_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21428\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48434\,
            ce => 'H',
            sr => \N__47862\
        );

    \pwm_generator_inst.threshold_4_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21464\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48434\,
            ce => 'H',
            sr => \N__47862\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100011011"
        )
    port map (
            in0 => \N__21253\,
            in1 => \N__21407\,
            in2 => \N__21348\,
            in3 => \N__20978\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48425\,
            ce => 'H',
            sr => \N__47869\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__21404\,
            in1 => \N__20963\,
            in2 => \N__21346\,
            in3 => \N__21254\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48425\,
            ce => 'H',
            sr => \N__47869\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__21252\,
            in1 => \N__21406\,
            in2 => \N__21347\,
            in3 => \N__21503\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48425\,
            ce => 'H',
            sr => \N__47869\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110101"
        )
    port map (
            in0 => \N__21405\,
            in1 => \N__21330\,
            in2 => \N__21273\,
            in3 => \N__21488\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48425\,
            ce => 'H',
            sr => \N__47869\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__21410\,
            in1 => \N__21289\,
            in2 => \N__21359\,
            in3 => \N__21470\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48413\,
            ce => 'H',
            sr => \N__47873\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__21409\,
            in1 => \N__21455\,
            in2 => \N__21358\,
            in3 => \N__21288\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48413\,
            ce => 'H',
            sr => \N__47873\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__21286\,
            in1 => \N__21355\,
            in2 => \N__21418\,
            in3 => \N__21449\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48413\,
            ce => 'H',
            sr => \N__47873\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__21287\,
            in1 => \N__21356\,
            in2 => \N__21419\,
            in3 => \N__21434\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48413\,
            ce => 'H',
            sr => \N__47873\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__21411\,
            in1 => \N__21357\,
            in2 => \N__21290\,
            in3 => \N__21116\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48406\,
            ce => 'H',
            sr => \N__47877\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21077\,
            in2 => \N__21110\,
            in3 => \N__21094\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21755\,
            in2 => \N__21800\,
            in3 => \N__21070\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21747\,
            in1 => \N__21731\,
            in2 => \N__21779\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21695\,
            in2 => \N__21725\,
            in3 => \N__21711\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21656\,
            in2 => \N__21689\,
            in3 => \N__21672\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21623\,
            in2 => \N__21650\,
            in3 => \N__21639\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21615\,
            in1 => \N__21590\,
            in2 => \N__21599\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21551\,
            in2 => \N__21584\,
            in3 => \N__21567\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21509\,
            in2 => \N__21545\,
            in3 => \N__21528\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21902\,
            in2 => \N__21938\,
            in3 => \N__21921\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21896\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48463\,
            ce => 'H',
            sr => \N__47824\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21962\,
            in1 => \N__21812\,
            in2 => \N__21956\,
            in3 => \N__22073\,
            lcout => \current_shift_inst.PI_CTRL.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22741\,
            in2 => \_gnd_net_\,
            in3 => \N__22363\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22721\,
            in1 => \N__22766\,
            in2 => \N__21815\,
            in3 => \N__22787\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_1_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21806\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48414\,
            ce => 'H',
            sr => \N__47863\
        );

    \pwm_generator_inst.threshold_2_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21788\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48414\,
            ce => 'H',
            sr => \N__47863\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21764\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27567\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24782\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => 'H',
            sr => \N__47817\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23516\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => 'H',
            sr => \N__47817\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27723\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28464\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22240\,
            in1 => \N__22255\,
            in2 => \N__22597\,
            in3 => \N__22270\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22559\,
            in1 => \N__22574\,
            in2 => \N__22601\,
            in3 => \N__22241\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22294\,
            in1 => \N__22256\,
            in2 => \N__22336\,
            in3 => \N__22271\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22537\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22519\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22573\,
            in1 => \N__22558\,
            in2 => \N__21947\,
            in3 => \N__21944\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22295\,
            in1 => \N__22745\,
            in2 => \N__22460\,
            in3 => \N__22364\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22831\,
            in2 => \_gnd_net_\,
            in3 => \N__22495\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22477\,
            in1 => \N__22802\,
            in2 => \N__22085\,
            in3 => \N__22817\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22801\,
            in2 => \_gnd_net_\,
            in3 => \N__22816\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22496\,
            in1 => \N__22520\,
            in2 => \N__22481\,
            in3 => \N__22541\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22459\,
            in1 => \N__22832\,
            in2 => \N__22082\,
            in3 => \N__22079\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22762\,
            in1 => \N__22786\,
            in2 => \N__22337\,
            in3 => \N__22720\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22067\,
            in1 => \N__22061\,
            in2 => \N__22052\,
            in3 => \N__22049\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21995\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48415\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_10_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__33524\,
            in1 => \N__23051\,
            in2 => \_gnd_net_\,
            in3 => \N__33141\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48380\,
            ce => 'H',
            sr => \N__47879\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22109\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22100\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__28298\,
            in1 => \N__28094\,
            in2 => \_gnd_net_\,
            in3 => \N__25196\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48453\,
            ce => 'H',
            sr => \N__47798\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31185\,
            in2 => \_gnd_net_\,
            in3 => \N__31601\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23704\,
            in2 => \_gnd_net_\,
            in3 => \N__24935\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__24965\,
            in1 => \N__24880\,
            in2 => \N__22091\,
            in3 => \N__27297\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110011"
        )
    port map (
            in0 => \N__23096\,
            in1 => \N__23656\,
            in2 => \N__22088\,
            in3 => \N__24745\,
            lcout => \current_shift_inst.PI_CTRL.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31600\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27406\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29696\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48435\,
            ce => 'H',
            sr => \N__47807\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29770\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48435\,
            ce => 'H',
            sr => \N__47807\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29860\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48435\,
            ce => 'H',
            sr => \N__47807\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27017\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48435\,
            ce => 'H',
            sr => \N__47807\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29818\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48435\,
            ce => 'H',
            sr => \N__47807\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23660\,
            in2 => \N__22226\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__48426\,
            ce => 'H',
            sr => \N__47812\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24934\,
            in2 => \N__23606\,
            in3 => \N__22160\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__48426\,
            ce => 'H',
            sr => \N__47812\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27302\,
            in2 => \N__23621\,
            in3 => \N__22139\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__48426\,
            ce => 'H',
            sr => \N__47812\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23705\,
            in2 => \N__23765\,
            in3 => \N__22112\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__48426\,
            ce => 'H',
            sr => \N__47812\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24976\,
            in2 => \N__22439\,
            in3 => \N__22412\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__48426\,
            ce => 'H',
            sr => \N__47812\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24886\,
            in2 => \N__22409\,
            in3 => \N__22376\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__48426\,
            ce => 'H',
            sr => \N__47812\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25024\,
            in2 => \N__22373\,
            in3 => \N__22340\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__48426\,
            ce => 'H',
            sr => \N__47812\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31919\,
            in2 => \N__24797\,
            in3 => \N__22307\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__48426\,
            ce => 'H',
            sr => \N__47812\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22304\,
            in2 => \N__31616\,
            in3 => \N__22274\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__48416\,
            ce => 'H',
            sr => \N__47818\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31267\,
            in2 => \N__29990\,
            in3 => \N__22259\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__48416\,
            ce => 'H',
            sr => \N__47818\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31189\,
            in2 => \N__29948\,
            in3 => \N__22244\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__48416\,
            ce => 'H',
            sr => \N__47818\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27402\,
            in2 => \N__23717\,
            in3 => \N__22229\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__48416\,
            ce => 'H',
            sr => \N__47818\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28471\,
            in2 => \N__28633\,
            in3 => \N__22577\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__48416\,
            ce => 'H',
            sr => \N__47818\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28602\,
            in2 => \N__27574\,
            in3 => \N__22562\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__48416\,
            ce => 'H',
            sr => \N__47818\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31740\,
            in2 => \N__28634\,
            in3 => \N__22544\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__48416\,
            ce => 'H',
            sr => \N__47818\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28606\,
            in2 => \N__31796\,
            in3 => \N__22523\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__48416\,
            ce => 'H',
            sr => \N__47818\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29516\,
            in2 => \N__28659\,
            in3 => \N__22499\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__48407\,
            ce => 'H',
            sr => \N__47825\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28638\,
            in2 => \N__31855\,
            in3 => \N__22484\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__48407\,
            ce => 'H',
            sr => \N__47825\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31685\,
            in2 => \N__28660\,
            in3 => \N__22463\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__48407\,
            ce => 'H',
            sr => \N__47825\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28642\,
            in2 => \N__27461\,
            in3 => \N__22442\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__48407\,
            ce => 'H',
            sr => \N__47825\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27724\,
            in2 => \N__28661\,
            in3 => \N__22820\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__48407\,
            ce => 'H',
            sr => \N__47825\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28646\,
            in2 => \N__27645\,
            in3 => \N__22805\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__48407\,
            ce => 'H',
            sr => \N__47825\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28725\,
            in2 => \N__28662\,
            in3 => \N__22790\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__48407\,
            ce => 'H',
            sr => \N__47825\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28650\,
            in2 => \N__27226\,
            in3 => \N__22769\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__48407\,
            ce => 'H',
            sr => \N__47825\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28397\,
            in2 => \N__28663\,
            in3 => \N__22748\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__48399\,
            ce => 'H',
            sr => \N__47834\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28654\,
            in2 => \N__28352\,
            in3 => \N__22724\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__48399\,
            ce => 'H',
            sr => \N__47834\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27772\,
            in2 => \N__28664\,
            in3 => \N__22706\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__48399\,
            ce => 'H',
            sr => \N__47834\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27903\,
            in1 => \N__28658\,
            in2 => \_gnd_net_\,
            in3 => \N__22703\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48399\,
            ce => 'H',
            sr => \N__47834\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22976\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22880\,
            in2 => \N__23162\,
            in3 => \N__23868\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22874\,
            in2 => \N__23327\,
            in3 => \N__23851\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22868\,
            in2 => \N__23150\,
            in3 => \N__23830\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22862\,
            in2 => \N__23315\,
            in3 => \N__23806\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22856\,
            in2 => \N__23303\,
            in3 => \N__23785\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22850\,
            in2 => \N__23189\,
            in3 => \N__24061\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24040\,
            in1 => \N__22844\,
            in2 => \N__23288\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24020\,
            in1 => \N__22838\,
            in2 => \N__23273\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22964\,
            in2 => \N__23177\,
            in3 => \N__23996\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23971\,
            in1 => \N__22940\,
            in2 => \N__22958\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22916\,
            in2 => \N__22934\,
            in3 => \N__23950\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22910\,
            in2 => \N__22991\,
            in3 => \N__23929\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22904\,
            in2 => \N__23234\,
            in3 => \N__23908\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22898\,
            in2 => \N__23264\,
            in3 => \N__24187\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22892\,
            in2 => \N__23336\,
            in3 => \N__24166\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22886\,
            in2 => \N__28859\,
            in3 => \N__25940\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23036\,
            in2 => \N__23015\,
            in3 => \N__24143\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24119\,
            in1 => \N__23030\,
            in2 => \N__23003\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23024\,
            in2 => \N__28874\,
            in3 => \N__24095\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23018\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25979\,
            in2 => \_gnd_net_\,
            in3 => \N__35601\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__30230\,
            in1 => \N__33992\,
            in2 => \_gnd_net_\,
            in3 => \N__34360\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48381\,
            ce => \N__28842\,
            sr => \N__47864\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34357\,
            in2 => \N__34010\,
            in3 => \N__30770\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48381\,
            ce => \N__28842\,
            sr => \N__47864\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34359\,
            in1 => \N__33743\,
            in2 => \N__34012\,
            in3 => \N__34177\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48381\,
            ce => \N__28842\,
            sr => \N__47864\
        );

    \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__34358\,
            in1 => \N__34176\,
            in2 => \N__34011\,
            in3 => \N__32569\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48381\,
            ce => \N__28842\,
            sr => \N__47864\
        );

    \delay_measurement_inst.delay_hc_reg_16_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__33514\,
            in1 => \N__23366\,
            in2 => \_gnd_net_\,
            in3 => \N__33142\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48376\,
            ce => 'H',
            sr => \N__47870\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25922\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48371\,
            ce => \N__24595\,
            sr => \N__47874\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25889\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48371\,
            ce => \N__24595\,
            sr => \N__47874\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__24391\,
            in1 => \N__24241\,
            in2 => \N__24521\,
            in3 => \N__29053\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_10_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33585\,
            in1 => \N__24392\,
            in2 => \_gnd_net_\,
            in3 => \N__33203\,
            lcout => \delay_measurement_inst.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI53F91_1_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24220\,
            in1 => \N__29052\,
            in2 => \_gnd_net_\,
            in3 => \N__26680\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__24242\,
            in1 => \N__30487\,
            in2 => \N__23039\,
            in3 => \N__24484\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_19_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33205\,
            in1 => \N__30285\,
            in2 => \_gnd_net_\,
            in3 => \N__24520\,
            lcout => \delay_measurement_inst.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_8_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24428\,
            in1 => \N__32659\,
            in2 => \_gnd_net_\,
            in3 => \N__33206\,
            lcout => \delay_measurement_inst.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_11_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33685\,
            in1 => \N__24368\,
            in2 => \_gnd_net_\,
            in3 => \N__33204\,
            lcout => \delay_measurement_inst.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__33452\,
            in1 => \N__23081\,
            in2 => \_gnd_net_\,
            in3 => \N__33132\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48359\,
            ce => 'H',
            sr => \N__47880\
        );

    \delay_measurement_inst.delay_hc_reg_11_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__33451\,
            in1 => \N__23075\,
            in2 => \_gnd_net_\,
            in3 => \N__33131\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48359\,
            ce => 'H',
            sr => \N__47880\
        );

    \delay_measurement_inst.delay_hc_reg_19_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__33138\,
            in1 => \N__33509\,
            in2 => \_gnd_net_\,
            in3 => \N__23069\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48353\,
            ce => 'H',
            sr => \N__47883\
        );

    \delay_measurement_inst.delay_hc_reg_12_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__33136\,
            in1 => \N__33507\,
            in2 => \_gnd_net_\,
            in3 => \N__23420\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48353\,
            ce => 'H',
            sr => \N__47883\
        );

    \delay_measurement_inst.delay_hc_reg_13_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__33137\,
            in1 => \N__33508\,
            in2 => \_gnd_net_\,
            in3 => \N__23441\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48353\,
            ce => 'H',
            sr => \N__47883\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23060\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__23541\,
            in1 => \N__38000\,
            in2 => \N__23575\,
            in3 => \N__23591\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48464\,
            ce => 'H',
            sr => \N__47788\
        );

    \phase_controller_inst2.state_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__35762\,
            in1 => \N__23543\,
            in2 => \N__23574\,
            in3 => \N__36818\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48454\,
            ce => 'H',
            sr => \N__47791\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111110011"
        )
    port map (
            in0 => \N__28301\,
            in1 => \N__27967\,
            in2 => \N__28132\,
            in3 => \N__25448\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48444\,
            ce => 'H',
            sr => \N__47795\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31739\,
            in1 => \N__25017\,
            in2 => \N__23222\,
            in3 => \N__23480\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23129\,
            in1 => \N__23105\,
            in2 => \N__23111\,
            in3 => \N__23138\,
            lcout => \current_shift_inst.PI_CTRL.N_74\,
            ltout => \current_shift_inst.PI_CTRL.N_74_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111110101"
        )
    port map (
            in0 => \N__27966\,
            in1 => \N__28302\,
            in2 => \N__23108\,
            in3 => \N__25409\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48444\,
            ce => 'H',
            sr => \N__47795\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36740\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36725\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36689\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29691\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30013\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31846\,
            in1 => \N__28396\,
            in2 => \N__27649\,
            in3 => \N__28729\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24778\,
            in1 => \N__23514\,
            in2 => \_gnd_net_\,
            in3 => \N__23743\,
            lcout => \current_shift_inst.PI_CTRL.un1_enablelt3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27219\,
            in1 => \N__27765\,
            in2 => \N__23090\,
            in3 => \N__23120\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24885\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24969\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27707\,
            in1 => \N__31678\,
            in2 => \N__31785\,
            in3 => \N__27885\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27641\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31774\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23698\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27442\,
            in1 => \N__28450\,
            in2 => \N__28351\,
            in3 => \N__31250\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28347\,
            in1 => \N__27443\,
            in2 => \N__27914\,
            in3 => \N__25009\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31249\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27550\,
            in1 => \N__27391\,
            in2 => \N__29503\,
            in3 => \N__31918\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI764B_28_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28392\,
            in2 => \_gnd_net_\,
            in3 => \N__31611\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_29_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23474\,
            in1 => \N__23210\,
            in2 => \N__30971\,
            in3 => \N__23204\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => \current_shift_inst.PI_CTRL.N_75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111110"
        )
    port map (
            in0 => \N__27886\,
            in1 => \N__28144\,
            in2 => \N__23192\,
            in3 => \N__25703\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48408\,
            ce => 'H',
            sr => \N__47813\
        );

    \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__34155\,
            in1 => \N__34004\,
            in2 => \N__30452\,
            in3 => \N__34340\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48400\,
            ce => \N__28831\,
            sr => \N__47819\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__34339\,
            in1 => \N__33643\,
            in2 => \N__34013\,
            in3 => \N__34156\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48400\,
            ce => \N__28831\,
            sr => \N__47819\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__34002\,
            in1 => \N__32875\,
            in2 => \_gnd_net_\,
            in3 => \N__32818\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48400\,
            ce => \N__28831\,
            sr => \N__47819\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__32819\,
            in1 => \N__34003\,
            in2 => \_gnd_net_\,
            in3 => \N__32795\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48400\,
            ce => \N__28831\,
            sr => \N__47819\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__35543\,
            in1 => \N__35425\,
            in2 => \N__35325\,
            in3 => \N__24029\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48395\,
            ce => 'H',
            sr => \N__47826\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__35424\,
            in1 => \N__35545\,
            in2 => \N__35324\,
            in3 => \N__24005\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48395\,
            ce => 'H',
            sr => \N__47826\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__35544\,
            in1 => \N__35426\,
            in2 => \N__35326\,
            in3 => \N__23981\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48395\,
            ce => 'H',
            sr => \N__47826\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__35542\,
            in1 => \N__35291\,
            in2 => \_gnd_net_\,
            in3 => \N__35423\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__35308\,
            in1 => \N__35431\,
            in2 => \N__35578\,
            in3 => \N__24128\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \N__47835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__35427\,
            in1 => \N__35546\,
            in2 => \N__35327\,
            in3 => \N__24104\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \N__47835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__35309\,
            in1 => \N__35432\,
            in2 => \N__35579\,
            in3 => \N__24077\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \N__47835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__35428\,
            in1 => \N__35547\,
            in2 => \N__35328\,
            in3 => \N__23840\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \N__47835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__35310\,
            in1 => \N__35433\,
            in2 => \N__35580\,
            in3 => \N__23819\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \N__47835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__35429\,
            in1 => \N__35548\,
            in2 => \N__35329\,
            in3 => \N__23795\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \N__47835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__35311\,
            in1 => \N__35434\,
            in2 => \N__35581\,
            in3 => \N__23774\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \N__47835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__35430\,
            in1 => \N__35549\,
            in2 => \N__35330\,
            in3 => \N__24050\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \N__47835\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__35301\,
            in1 => \N__23960\,
            in2 => \N__35584\,
            in3 => \N__35440\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48387\,
            ce => 'H',
            sr => \N__47843\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__25978\,
            in1 => \N__23872\,
            in2 => \_gnd_net_\,
            in3 => \N__35609\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__35304\,
            in1 => \N__35527\,
            in2 => \N__23237\,
            in3 => \N__35441\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48387\,
            ce => 'H',
            sr => \N__47843\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__35435\,
            in1 => \N__35305\,
            in2 => \N__35571\,
            in3 => \N__23939\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48387\,
            ce => 'H',
            sr => \N__47843\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__35302\,
            in1 => \N__35438\,
            in2 => \N__35582\,
            in3 => \N__23918\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48387\,
            ce => 'H',
            sr => \N__47843\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__35436\,
            in1 => \N__35306\,
            in2 => \N__35572\,
            in3 => \N__23897\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48387\,
            ce => 'H',
            sr => \N__47843\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__35303\,
            in1 => \N__35439\,
            in2 => \N__35583\,
            in3 => \N__24176\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48387\,
            ce => 'H',
            sr => \N__47843\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__35437\,
            in1 => \N__35307\,
            in2 => \N__35573\,
            in3 => \N__24155\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48387\,
            ce => 'H',
            sr => \N__47843\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__33945\,
            in1 => \N__34341\,
            in2 => \N__34506\,
            in3 => \N__34097\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48382\,
            ce => \N__28832\,
            sr => \N__47851\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34099\,
            in1 => \N__34424\,
            in2 => \N__34362\,
            in3 => \N__33956\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48382\,
            ce => \N__28832\,
            sr => \N__47851\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33946\,
            in1 => \N__34100\,
            in2 => \N__34058\,
            in3 => \N__34356\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48382\,
            ce => \N__28832\,
            sr => \N__47851\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34101\,
            in1 => \N__33947\,
            in2 => \N__34363\,
            in3 => \N__32431\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48382\,
            ce => \N__28832\,
            sr => \N__47851\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32369\,
            in1 => \N__34342\,
            in2 => \N__33985\,
            in3 => \N__34102\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48382\,
            ce => \N__28832\,
            sr => \N__47851\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34103\,
            in1 => \N__33948\,
            in2 => \N__34364\,
            in3 => \N__32724\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48382\,
            ce => \N__28832\,
            sr => \N__47851\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32670\,
            in1 => \N__34343\,
            in2 => \N__33986\,
            in3 => \N__34104\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48382\,
            ce => \N__28832\,
            sr => \N__47851\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__34098\,
            in1 => \N__30362\,
            in2 => \N__34361\,
            in3 => \N__33955\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48382\,
            ce => \N__28832\,
            sr => \N__47851\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__33140\,
            in1 => \N__23372\,
            in2 => \N__33523\,
            in3 => \_gnd_net_\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48377\,
            ce => 'H',
            sr => \N__47858\
        );

    \phase_controller_inst2.S2_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23579\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48377\,
            ce => 'H',
            sr => \N__47858\
        );

    \delay_measurement_inst.delay_hc_reg_17_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__24254\,
            in1 => \N__33500\,
            in2 => \_gnd_net_\,
            in3 => \N__33139\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48377\,
            ce => 'H',
            sr => \N__47858\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_7_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33273\,
            in1 => \N__32723\,
            in2 => \_gnd_net_\,
            in3 => \N__24450\,
            lcout => \delay_measurement_inst.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__24414\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24449\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_16_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__33272\,
            in1 => \_gnd_net_\,
            in2 => \N__32920\,
            in3 => \N__24571\,
            lcout => \delay_measurement_inst.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_14_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30349\,
            in1 => \N__24287\,
            in2 => \_gnd_net_\,
            in3 => \N__33271\,
            lcout => \delay_measurement_inst.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24304\,
            in1 => \N__24361\,
            in2 => \N__24337\,
            in3 => \N__24385\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFRS4_9_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010000"
        )
    port map (
            in0 => \N__28758\,
            in1 => \N__23360\,
            in2 => \N__23354\,
            in3 => \N__23351\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24303\,
            in1 => \N__28757\,
            in2 => \N__24572\,
            in3 => \N__24471\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24546\,
            in1 => \N__24516\,
            in2 => \N__28977\,
            in3 => \N__24570\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JGD6_14_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__26764\,
            in1 => \N__24286\,
            in2 => \N__23345\,
            in3 => \N__23342\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_6_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24472\,
            in1 => \N__24415\,
            in2 => \_gnd_net_\,
            in3 => \N__24451\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000100"
        )
    port map (
            in0 => \N__23414\,
            in1 => \N__24285\,
            in2 => \N__23408\,
            in3 => \N__28759\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_4_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24219\,
            in1 => \N__32426\,
            in2 => \_gnd_net_\,
            in3 => \N__33202\,
            lcout => \delay_measurement_inst.N_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24284\,
            in1 => \N__24360\,
            in2 => \N__24336\,
            in3 => \N__26762\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJAU73_7_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24427\,
            in1 => \N__24455\,
            in2 => \N__23405\,
            in3 => \N__23402\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_17_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__29018\,
            in1 => \N__23450\,
            in2 => \N__23396\,
            in3 => \N__24698\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__26763\,
            in1 => \N__23393\,
            in2 => \N__23384\,
            in3 => \N__23381\,
            lcout => \delay_measurement_inst.un1_elapsed_time_hc\,
            ltout => \delay_measurement_inst.un1_elapsed_time_hc_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_3_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32790\,
            in2 => \N__23375\,
            in3 => \N__24240\,
            lcout => \delay_measurement_inst.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__24221\,
            in1 => \_gnd_net_\,
            in2 => \N__30486\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_17_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24550\,
            in1 => \N__28981\,
            in2 => \N__23462\,
            in3 => \N__23459\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30422\,
            in1 => \N__24485\,
            in2 => \_gnd_net_\,
            in3 => \N__33259\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.N_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_6_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110101"
        )
    port map (
            in0 => \N__33130\,
            in1 => \_gnd_net_\,
            in2 => \N__23444\,
            in3 => \N__33378\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48354\,
            ce => 'H',
            sr => \N__47878\
        );

    \delay_measurement_inst.delay_hc_reg_25_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__33377\,
            in1 => \N__33260\,
            in2 => \N__29207\,
            in3 => \N__33129\,
            lcout => measured_delay_hc_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48354\,
            ce => 'H',
            sr => \N__47878\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_13_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34466\,
            in1 => \N__24308\,
            in2 => \_gnd_net_\,
            in3 => \N__33262\,
            lcout => \delay_measurement_inst.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29237\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29271\,
            in2 => \_gnd_net_\,
            in3 => \N__29236\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_302_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_12_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33728\,
            in1 => \N__24341\,
            in2 => \_gnd_net_\,
            in3 => \N__33261\,
            lcout => \delay_measurement_inst.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_state_0_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__24815\,
            in1 => \N__24831\,
            in2 => \_gnd_net_\,
            in3 => \N__30563\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48465\,
            ce => \N__35904\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__24814\,
            in1 => \N__24832\,
            in2 => \N__47927\,
            in3 => \N__30569\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48455\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37996\,
            in2 => \_gnd_net_\,
            in3 => \N__23590\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27560\,
            in1 => \N__27401\,
            in2 => \N__29522\,
            in3 => \N__31912\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23564\,
            in2 => \_gnd_net_\,
            in3 => \N__23542\,
            lcout => \phase_controller_inst2.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__31512\,
            in1 => \N__29819\,
            in2 => \N__23515\,
            in3 => \N__26966\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23507\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23702\,
            in1 => \N__27301\,
            in2 => \N__24884\,
            in3 => \N__24925\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__24964\,
            in1 => \N__23648\,
            in2 => \N__23483\,
            in3 => \N__24728\,
            lcout => \current_shift_inst.PI_CTRL.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28463\,
            in1 => \N__31177\,
            in2 => \N__27776\,
            in3 => \N__31260\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23742\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25016\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__31517\,
            in1 => \N__29692\,
            in2 => \N__23655\,
            in3 => \N__27113\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23644\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__27915\,
            in1 => \N__28282\,
            in2 => \N__28130\,
            in3 => \N__25100\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48427\,
            ce => 'H',
            sr => \N__47796\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__28279\,
            in1 => \N__28084\,
            in2 => \N__27965\,
            in3 => \N__25352\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48427\,
            ce => 'H',
            sr => \N__47796\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111110"
        )
    port map (
            in0 => \N__28083\,
            in1 => \N__28280\,
            in2 => \N__27964\,
            in3 => \N__25325\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48427\,
            ce => 'H',
            sr => \N__47796\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111101010100"
        )
    port map (
            in0 => \N__25283\,
            in1 => \N__28281\,
            in2 => \N__28131\,
            in3 => \N__27922\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48427\,
            ce => 'H',
            sr => \N__47796\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29906\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48417\,
            ce => 'H',
            sr => \N__47799\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29933\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48417\,
            ce => 'H',
            sr => \N__47799\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011111110"
        )
    port map (
            in0 => \N__28122\,
            in1 => \N__27971\,
            in2 => \N__28304\,
            in3 => \N__25730\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48417\,
            ce => 'H',
            sr => \N__47799\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000111"
        )
    port map (
            in0 => \N__25070\,
            in1 => \N__28285\,
            in2 => \N__28000\,
            in3 => \N__28125\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48417\,
            ce => 'H',
            sr => \N__47799\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011111110"
        )
    port map (
            in0 => \N__28121\,
            in1 => \N__27970\,
            in2 => \N__28303\,
            in3 => \N__25370\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48417\,
            ce => 'H',
            sr => \N__47799\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110101110"
        )
    port map (
            in0 => \N__27969\,
            in1 => \N__28284\,
            in2 => \N__25580\,
            in3 => \N__28124\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48417\,
            ce => 'H',
            sr => \N__47799\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110101110"
        )
    port map (
            in0 => \N__27968\,
            in1 => \N__28283\,
            in2 => \N__25295\,
            in3 => \N__28123\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48417\,
            ce => 'H',
            sr => \N__47799\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__31469\,
            in1 => \N__30043\,
            in2 => \N__23703\,
            in3 => \N__27080\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111001111"
        )
    port map (
            in0 => \N__28251\,
            in1 => \N__28129\,
            in2 => \N__28003\,
            in3 => \N__25037\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48409\,
            ce => 'H',
            sr => \N__47803\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__28249\,
            in1 => \N__28127\,
            in2 => \N__28001\,
            in3 => \N__25607\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48409\,
            ce => 'H',
            sr => \N__47803\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__28250\,
            in1 => \N__28128\,
            in2 => \N__28002\,
            in3 => \N__25550\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48409\,
            ce => 'H',
            sr => \N__47803\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101001110"
        )
    port map (
            in0 => \N__28126\,
            in1 => \N__27981\,
            in2 => \N__25526\,
            in3 => \N__28252\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48409\,
            ce => 'H',
            sr => \N__47803\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29885\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__47808\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101001110"
        )
    port map (
            in0 => \N__28147\,
            in1 => \N__27985\,
            in2 => \N__25640\,
            in3 => \N__28247\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__47808\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__25229\,
            in1 => \_gnd_net_\,
            in2 => \N__28292\,
            in3 => \N__28152\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__47808\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101001110"
        )
    port map (
            in0 => \N__28148\,
            in1 => \N__27986\,
            in2 => \N__25514\,
            in3 => \N__28248\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__47808\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__28241\,
            in1 => \N__28150\,
            in2 => \N__28004\,
            in3 => \N__25499\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__47808\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101001110"
        )
    port map (
            in0 => \N__28149\,
            in1 => \N__27987\,
            in2 => \N__25490\,
            in3 => \N__28246\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__47808\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__28242\,
            in1 => \N__28151\,
            in2 => \N__28005\,
            in3 => \N__25478\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__47808\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30047\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \N__47808\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27716\,
            in1 => \N__28712\,
            in2 => \N__27218\,
            in3 => \N__27629\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__28253\,
            in1 => \N__28145\,
            in2 => \N__28006\,
            in3 => \N__25679\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48396\,
            ce => 'H',
            sr => \N__47814\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28711\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__28254\,
            in1 => \N__28146\,
            in2 => \N__28007\,
            in3 => \N__25661\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48396\,
            ce => 'H',
            sr => \N__47814\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27208\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23888\,
            in2 => \N__23876\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23852\,
            in2 => \_gnd_net_\,
            in3 => \N__23834\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23831\,
            in2 => \N__25760\,
            in3 => \N__23813\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23810\,
            in3 => \N__23789\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23786\,
            in2 => \_gnd_net_\,
            in3 => \N__23768\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24062\,
            in2 => \_gnd_net_\,
            in3 => \N__24044\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24041\,
            in2 => \_gnd_net_\,
            in3 => \N__24023\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24019\,
            in2 => \_gnd_net_\,
            in3 => \N__23999\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23995\,
            in2 => \_gnd_net_\,
            in3 => \N__23975\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23972\,
            in2 => \_gnd_net_\,
            in3 => \N__23954\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23951\,
            in2 => \_gnd_net_\,
            in3 => \N__23933\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23930\,
            in2 => \_gnd_net_\,
            in3 => \N__23912\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23909\,
            in2 => \_gnd_net_\,
            in3 => \N__23891\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24188\,
            in2 => \_gnd_net_\,
            in3 => \N__24170\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24167\,
            in2 => \_gnd_net_\,
            in3 => \N__24149\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25939\,
            in2 => \_gnd_net_\,
            in3 => \N__24146\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24142\,
            in2 => \_gnd_net_\,
            in3 => \N__24122\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24118\,
            in2 => \_gnd_net_\,
            in3 => \N__24098\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24094\,
            in2 => \_gnd_net_\,
            in3 => \N__24080\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30765\,
            in1 => \N__32927\,
            in2 => \N__30296\,
            in3 => \N__30238\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__34429\,
            in1 => \N__30357\,
            in2 => \N__24071\,
            in3 => \N__24260\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt30\,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlt30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto31_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36206\,
            in2 => \N__24266\,
            in3 => \N__34303\,
            lcout => \phase_controller_inst1.stoper_hc.un1_start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33750\,
            in1 => \N__33698\,
            in2 => \N__34502\,
            in3 => \N__33581\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010000"
        )
    port map (
            in0 => \N__33635\,
            in1 => \N__24248\,
            in2 => \N__24263\,
            in3 => \N__30314\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_ibuf_gb_io_RNI79U7_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47922\,
            lcout => red_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_17_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30229\,
            in1 => \N__24551\,
            in2 => \_gnd_net_\,
            in3 => \N__33289\,
            lcout => \delay_measurement_inst.N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32666\,
            in2 => \_gnd_net_\,
            in3 => \N__32716\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25855\,
            in2 => \N__25921\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__48366\,
            ce => \N__24599\,
            sr => \N__47859\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25882\,
            in2 => \N__25832\,
            in3 => \N__24194\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__48366\,
            ce => \N__24599\,
            sr => \N__47859\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25856\,
            in2 => \N__26194\,
            in3 => \N__24191\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__48366\,
            ce => \N__24599\,
            sr => \N__47859\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25828\,
            in2 => \N__26164\,
            in3 => \N__24458\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__48366\,
            ce => \N__24599\,
            sr => \N__47859\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26137\,
            in2 => \N__26195\,
            in3 => \N__24431\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__48366\,
            ce => \N__24599\,
            sr => \N__47859\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26116\,
            in2 => \N__26165\,
            in3 => \N__24398\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__48366\,
            ce => \N__24599\,
            sr => \N__47859\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26138\,
            in2 => \N__26089\,
            in3 => \N__24395\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__48366\,
            ce => \N__24599\,
            sr => \N__47859\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26117\,
            in2 => \N__26056\,
            in3 => \N__24371\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__48366\,
            ce => \N__24599\,
            sr => \N__47859\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26093\,
            in2 => \N__26029\,
            in3 => \N__24344\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__48360\,
            ce => \N__24598\,
            sr => \N__47865\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26002\,
            in2 => \N__26063\,
            in3 => \N__24311\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__48360\,
            ce => \N__24598\,
            sr => \N__47865\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26428\,
            in2 => \N__26030\,
            in3 => \N__24290\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__48360\,
            ce => \N__24598\,
            sr => \N__47865\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26003\,
            in2 => \N__26407\,
            in3 => \N__24578\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__48360\,
            ce => \N__24598\,
            sr => \N__47865\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26429\,
            in2 => \N__26381\,
            in3 => \N__24575\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__48360\,
            ce => \N__24598\,
            sr => \N__47865\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26350\,
            in2 => \N__26408\,
            in3 => \N__24554\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__48360\,
            ce => \N__24598\,
            sr => \N__47865\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26377\,
            in2 => \N__26326\,
            in3 => \N__24527\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__48360\,
            ce => \N__24598\,
            sr => \N__47865\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26351\,
            in2 => \N__26290\,
            in3 => \N__24524\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__48360\,
            ce => \N__24598\,
            sr => \N__47865\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26327\,
            in2 => \N__26263\,
            in3 => \N__24497\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__48355\,
            ce => \N__24597\,
            sr => \N__47871\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26236\,
            in2 => \N__26297\,
            in3 => \N__24494\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__48355\,
            ce => \N__24597\,
            sr => \N__47871\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26215\,
            in2 => \N__26264\,
            in3 => \N__24491\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__48355\,
            ce => \N__24597\,
            sr => \N__47871\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26237\,
            in2 => \N__26641\,
            in3 => \N__24488\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__48355\,
            ce => \N__24597\,
            sr => \N__47871\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26216\,
            in2 => \N__26615\,
            in3 => \N__24626\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__48355\,
            ce => \N__24597\,
            sr => \N__47871\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26584\,
            in2 => \N__26642\,
            in3 => \N__24623\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__48355\,
            ce => \N__24597\,
            sr => \N__47871\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26611\,
            in2 => \N__26557\,
            in3 => \N__24620\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__48355\,
            ce => \N__24597\,
            sr => \N__47871\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26585\,
            in2 => \N__26524\,
            in3 => \N__24617\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__48355\,
            ce => \N__24597\,
            sr => \N__47871\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26494\,
            in2 => \N__26561\,
            in3 => \N__24614\,
            lcout => \delay_measurement_inst.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__48349\,
            ce => \N__24596\,
            sr => \N__47875\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26467\,
            in2 => \N__26531\,
            in3 => \N__24611\,
            lcout => \delay_measurement_inst.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__48349\,
            ce => \N__24596\,
            sr => \N__47875\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26447\,
            in2 => \N__26498\,
            in3 => \N__24608\,
            lcout => \delay_measurement_inst.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__48349\,
            ce => \N__24596\,
            sr => \N__47875\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26468\,
            in2 => \N__26783\,
            in3 => \N__24605\,
            lcout => \delay_measurement_inst.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__48349\,
            ce => \N__24596\,
            sr => \N__47875\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24602\,
            lcout => \delay_measurement_inst.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48349\,
            ce => \N__24596\,
            sr => \N__47875\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26668\,
            in1 => \N__24688\,
            in2 => \N__29119\,
            in3 => \N__30640\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUV512_20_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__29035\,
            in1 => \N__33376\,
            in2 => \N__24701\,
            in3 => \N__26702\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_28_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29137\,
            in1 => \N__24689\,
            in2 => \_gnd_net_\,
            in3 => \N__33316\,
            lcout => \delay_measurement_inst.N_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_28_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__24680\,
            in1 => \N__33437\,
            in2 => \_gnd_net_\,
            in3 => \N__33143\,
            lcout => measured_delay_hc_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48340\,
            ce => 'H',
            sr => \N__47881\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24656\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24644\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48446\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43419\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24632\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48446\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__24813\,
            in1 => \N__24833\,
            in2 => \_gnd_net_\,
            in3 => \N__30564\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48437\,
            ce => 'H',
            sr => \N__47774\
        );

    \delay_measurement_inst.prev_hc_sig_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.prev_hc_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48437\,
            ce => 'H',
            sr => \N__47774\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36013\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48429\,
            ce => 'H',
            sr => \N__47778\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29740\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48429\,
            ce => 'H',
            sr => \N__47778\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__31521\,
            in1 => \N__29771\,
            in2 => \N__24771\,
            in3 => \N__27140\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24761\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__28299\,
            in1 => \N__28101\,
            in2 => \_gnd_net_\,
            in3 => \N__25160\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48419\,
            ce => 'H',
            sr => \N__47784\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__28300\,
            in1 => \N__28102\,
            in2 => \_gnd_net_\,
            in3 => \N__25127\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48419\,
            ce => 'H',
            sr => \N__47784\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24727\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__27131\,
            in1 => \N__29741\,
            in2 => \N__24744\,
            in3 => \N__31522\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__26975\,
            in1 => \N__29861\,
            in2 => \N__25256\,
            in3 => \N__31514\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__31547\,
            in1 => \N__31519\,
            in2 => \N__25028\,
            in3 => \N__27044\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31513\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__29651\,
            in1 => \N__31520\,
            in2 => \N__31916\,
            in3 => \N__27170\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011111111"
        )
    port map (
            in0 => \N__27065\,
            in1 => \N__29609\,
            in2 => \N__24980\,
            in3 => \N__31516\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__31515\,
            in1 => \N__30014\,
            in2 => \N__24933\,
            in3 => \N__27092\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31735\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__29630\,
            in1 => \N__31518\,
            in2 => \N__24893\,
            in3 => \N__27053\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24844\,
            in2 => \N__24848\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25252\,
            in2 => \N__25238\,
            in3 => \N__25220\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25217\,
            in2 => \N__25208\,
            in3 => \N__25184\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25181\,
            in2 => \N__25172\,
            in3 => \N__25151\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25148\,
            in2 => \N__25139\,
            in3 => \N__25118\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25115\,
            in2 => \N__25109\,
            in3 => \N__25094\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25091\,
            in2 => \N__25085\,
            in3 => \N__25061\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25769\,
            in2 => \N__27323\,
            in3 => \N__25058\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25055\,
            in2 => \N__25049\,
            in3 => \N__25031\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \bfn_10_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25472\,
            in2 => \N__25463\,
            in3 => \N__25436\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25433\,
            in2 => \N__25424\,
            in3 => \N__25397\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25394\,
            in2 => \N__25385\,
            in3 => \N__25364\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25361\,
            in2 => \N__31868\,
            in3 => \N__25343\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31556\,
            in2 => \N__25340\,
            in3 => \N__25313\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31217\,
            in2 => \N__25310\,
            in3 => \N__25286\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31133\,
            in2 => \N__29666\,
            in3 => \N__25274\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27350\,
            in2 => \N__25271\,
            in3 => \N__25628\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28412\,
            in2 => \N__25625\,
            in3 => \N__25601\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27509\,
            in2 => \N__25598\,
            in3 => \N__25568\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29540\,
            in2 => \N__25565\,
            in3 => \N__25544\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27467\,
            in2 => \N__25541\,
            in3 => \N__25517\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27485\,
            in2 => \N__29465\,
            in3 => \N__25502\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27338\,
            in2 => \N__26954\,
            in3 => \N__25493\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27497\,
            in2 => \N__30953\,
            in3 => \N__25481\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27413\,
            in2 => \N__25799\,
            in3 => \N__25751\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27671\,
            in2 => \N__25748\,
            in3 => \N__25721\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27596\,
            in2 => \N__25718\,
            in3 => \N__25691\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28688\,
            in2 => \N__25688\,
            in3 => \N__25673\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27182\,
            in2 => \N__25670\,
            in3 => \N__25655\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25790\,
            in2 => \N__28681\,
            in3 => \N__25652\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28677\,
            in2 => \N__25778\,
            in3 => \N__25649\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25784\,
            in2 => \N__28682\,
            in3 => \N__25646\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27879\,
            in1 => \N__31523\,
            in2 => \_gnd_net_\,
            in3 => \N__25643\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27453\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28374\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27747\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28326\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27275\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25974\,
            in2 => \_gnd_net_\,
            in3 => \N__35619\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__35502\,
            in1 => \N__35289\,
            in2 => \_gnd_net_\,
            in3 => \N__35377\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__45523\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45482\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34612\,
            in2 => \_gnd_net_\,
            in3 => \N__33798\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__35491\,
            in1 => \N__28880\,
            in2 => \N__25982\,
            in3 => \N__45488\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48372\,
            ce => 'H',
            sr => \N__47820\
        );

    \phase_controller_inst1.state_2_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__33799\,
            in1 => \N__30703\,
            in2 => \N__34616\,
            in3 => \N__30678\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48372\,
            ce => 'H',
            sr => \N__47820\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35288\,
            in2 => \_gnd_net_\,
            in3 => \N__35376\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed11\,
            ltout => \phase_controller_inst1.stoper_hc.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011011000"
        )
    port map (
            in0 => \N__25955\,
            in1 => \N__30679\,
            in2 => \N__25949\,
            in3 => \N__35631\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48372\,
            ce => 'H',
            sr => \N__47820\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__35290\,
            in1 => \N__35492\,
            in2 => \N__35422\,
            in3 => \N__25946\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48372\,
            ce => 'H',
            sr => \N__47820\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26936\,
            in1 => \N__25908\,
            in2 => \_gnd_net_\,
            in3 => \N__25892\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__48367\,
            ce => \N__28948\,
            sr => \N__47827\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26932\,
            in1 => \N__25875\,
            in2 => \_gnd_net_\,
            in3 => \N__25859\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__48367\,
            ce => \N__28948\,
            sr => \N__47827\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26937\,
            in1 => \N__25854\,
            in2 => \_gnd_net_\,
            in3 => \N__25835\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__48367\,
            ce => \N__28948\,
            sr => \N__47827\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26933\,
            in1 => \N__25824\,
            in2 => \_gnd_net_\,
            in3 => \N__25802\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__48367\,
            ce => \N__28948\,
            sr => \N__47827\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26938\,
            in1 => \N__26182\,
            in2 => \_gnd_net_\,
            in3 => \N__26168\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__48367\,
            ce => \N__28948\,
            sr => \N__47827\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26934\,
            in1 => \N__26157\,
            in2 => \_gnd_net_\,
            in3 => \N__26141\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__48367\,
            ce => \N__28948\,
            sr => \N__47827\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26939\,
            in1 => \N__26136\,
            in2 => \_gnd_net_\,
            in3 => \N__26120\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__48367\,
            ce => \N__28948\,
            sr => \N__47827\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26935\,
            in1 => \N__26110\,
            in2 => \_gnd_net_\,
            in3 => \N__26096\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__48367\,
            ce => \N__28948\,
            sr => \N__47827\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26927\,
            in1 => \N__26085\,
            in2 => \_gnd_net_\,
            in3 => \N__26066\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__48362\,
            ce => \N__28949\,
            sr => \N__47836\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26931\,
            in1 => \N__26055\,
            in2 => \_gnd_net_\,
            in3 => \N__26033\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__48362\,
            ce => \N__28949\,
            sr => \N__47836\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26924\,
            in1 => \N__26022\,
            in2 => \_gnd_net_\,
            in3 => \N__26006\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__48362\,
            ce => \N__28949\,
            sr => \N__47836\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26928\,
            in1 => \N__26001\,
            in2 => \_gnd_net_\,
            in3 => \N__25985\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__48362\,
            ce => \N__28949\,
            sr => \N__47836\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26925\,
            in1 => \N__26427\,
            in2 => \_gnd_net_\,
            in3 => \N__26411\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__48362\,
            ce => \N__28949\,
            sr => \N__47836\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26929\,
            in1 => \N__26400\,
            in2 => \_gnd_net_\,
            in3 => \N__26384\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__48362\,
            ce => \N__28949\,
            sr => \N__47836\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26926\,
            in1 => \N__26373\,
            in2 => \_gnd_net_\,
            in3 => \N__26354\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__48362\,
            ce => \N__28949\,
            sr => \N__47836\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26930\,
            in1 => \N__26344\,
            in2 => \_gnd_net_\,
            in3 => \N__26330\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__48362\,
            ce => \N__28949\,
            sr => \N__47836\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26910\,
            in1 => \N__26322\,
            in2 => \_gnd_net_\,
            in3 => \N__26300\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__48356\,
            ce => \N__28940\,
            sr => \N__47847\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26917\,
            in1 => \N__26289\,
            in2 => \_gnd_net_\,
            in3 => \N__26267\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__48356\,
            ce => \N__28940\,
            sr => \N__47847\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26911\,
            in1 => \N__26256\,
            in2 => \_gnd_net_\,
            in3 => \N__26240\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__48356\,
            ce => \N__28940\,
            sr => \N__47847\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26914\,
            in1 => \N__26235\,
            in2 => \_gnd_net_\,
            in3 => \N__26219\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__48356\,
            ce => \N__28940\,
            sr => \N__47847\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26912\,
            in1 => \N__26214\,
            in2 => \_gnd_net_\,
            in3 => \N__26198\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__48356\,
            ce => \N__28940\,
            sr => \N__47847\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26915\,
            in1 => \N__26634\,
            in2 => \_gnd_net_\,
            in3 => \N__26618\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__48356\,
            ce => \N__28940\,
            sr => \N__47847\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26913\,
            in1 => \N__26607\,
            in2 => \_gnd_net_\,
            in3 => \N__26588\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__48356\,
            ce => \N__28940\,
            sr => \N__47847\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26916\,
            in1 => \N__26578\,
            in2 => \_gnd_net_\,
            in3 => \N__26564\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__48356\,
            ce => \N__28940\,
            sr => \N__47847\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26918\,
            in1 => \N__26553\,
            in2 => \_gnd_net_\,
            in3 => \N__26534\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__48350\,
            ce => \N__28944\,
            sr => \N__47852\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26922\,
            in1 => \N__26523\,
            in2 => \_gnd_net_\,
            in3 => \N__26501\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__48350\,
            ce => \N__28944\,
            sr => \N__47852\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26919\,
            in1 => \N__26487\,
            in2 => \_gnd_net_\,
            in3 => \N__26471\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__48350\,
            ce => \N__28944\,
            sr => \N__47852\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26923\,
            in1 => \N__26466\,
            in2 => \_gnd_net_\,
            in3 => \N__26450\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__48350\,
            ce => \N__28944\,
            sr => \N__47852\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26920\,
            in1 => \N__26446\,
            in2 => \_gnd_net_\,
            in3 => \N__26432\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__48350\,
            ce => \N__28944\,
            sr => \N__47852\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__26779\,
            in1 => \N__26921\,
            in2 => \_gnd_net_\,
            in3 => \N__26786\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48350\,
            ce => \N__28944\,
            sr => \N__47852\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_15_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34400\,
            in1 => \N__26765\,
            in2 => \_gnd_net_\,
            in3 => \N__33293\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.N_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_15_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33414\,
            in2 => \N__26744\,
            in3 => \N__33077\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48346\,
            ce => 'H',
            sr => \N__47860\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26741\,
            in1 => \N__26735\,
            in2 => \N__26729\,
            in3 => \N__26720\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26714\,
            in2 => \_gnd_net_\,
            in3 => \N__26708\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI45SG1_21_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26696\,
            in3 => \N__26693\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_1_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32866\,
            in1 => \N__33315\,
            in2 => \_gnd_net_\,
            in3 => \N__26687\,
            lcout => \delay_measurement_inst.N_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_27_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26669\,
            in1 => \N__29096\,
            in2 => \_gnd_net_\,
            in3 => \N__33317\,
            lcout => \delay_measurement_inst.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35831\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48330\,
            ce => 'H',
            sr => \N__47884\
        );

    \delay_measurement_inst.tr_state_0_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__29366\,
            in1 => \N__29343\,
            in2 => \_gnd_net_\,
            in3 => \N__29327\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48458\,
            ce => \N__35927\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__39072\,
            in1 => \N__39114\,
            in2 => \N__38748\,
            in3 => \N__42747\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__41433\,
            in1 => \N__41288\,
            in2 => \_gnd_net_\,
            in3 => \N__37276\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48438\,
            ce => \N__30869\,
            sr => \N__47765\
        );

    \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__29414\,
            in1 => \N__41429\,
            in2 => \_gnd_net_\,
            in3 => \N__40985\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48438\,
            ce => \N__30869\,
            sr => \N__47765\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__40880\,
            in1 => \_gnd_net_\,
            in2 => \N__41435\,
            in3 => \N__37275\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48438\,
            ce => \N__30869\,
            sr => \N__47765\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__37277\,
            in1 => \N__41434\,
            in2 => \_gnd_net_\,
            in3 => \N__41234\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48438\,
            ce => \N__30869\,
            sr => \N__47765\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31854\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39063\,
            in1 => \N__39113\,
            in2 => \N__38747\,
            in3 => \N__42746\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__40936\,
            in1 => \N__41128\,
            in2 => \N__30890\,
            in3 => \N__37261\,
            lcout => \delay_measurement_inst.N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101110"
        )
    port map (
            in0 => \N__37262\,
            in1 => \N__40937\,
            in2 => \N__40835\,
            in3 => \N__40984\,
            lcout => \delay_measurement_inst.N_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__37582\,
            in1 => \N__45487\,
            in2 => \N__28789\,
            in3 => \N__27038\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48420\,
            ce => 'H',
            sr => \N__47775\
        );

    \phase_controller_inst1.start_timer_tr_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__45486\,
            in1 => \N__43601\,
            in2 => \N__27029\,
            in3 => \N__43855\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48420\,
            ce => 'H',
            sr => \N__47775\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26999\,
            in2 => \_gnd_net_\,
            in3 => \N__27010\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26993\,
            in2 => \_gnd_net_\,
            in3 => \N__29932\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26987\,
            in2 => \_gnd_net_\,
            in3 => \N__29905\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26981\,
            in2 => \_gnd_net_\,
            in3 => \N__29881\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29588\,
            in2 => \_gnd_net_\,
            in3 => \N__26969\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29432\,
            in2 => \_gnd_net_\,
            in3 => \N__26957\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29582\,
            in2 => \_gnd_net_\,
            in3 => \N__27134\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29426\,
            in2 => \_gnd_net_\,
            in3 => \N__27125\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27122\,
            in2 => \_gnd_net_\,
            in3 => \N__27104\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_8\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27101\,
            in2 => \_gnd_net_\,
            in3 => \N__27086\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29447\,
            in3 => \N__27083\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29438\,
            in2 => \_gnd_net_\,
            in3 => \N__27068\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29604\,
            in2 => \_gnd_net_\,
            in3 => \N__27056\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29625\,
            in2 => \_gnd_net_\,
            in3 => \N__27047\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31546\,
            in2 => \_gnd_net_\,
            in3 => \N__27173\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29646\,
            in2 => \_gnd_net_\,
            in3 => \N__27164\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31634\,
            in2 => \_gnd_net_\,
            in3 => \N__27161\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31298\,
            in2 => \_gnd_net_\,
            in3 => \N__27158\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31205\,
            in2 => \_gnd_net_\,
            in3 => \N__27155\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31117\,
            in2 => \_gnd_net_\,
            in3 => \N__27152\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31063\,
            in2 => \_gnd_net_\,
            in3 => \N__27149\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28574\,
            in2 => \_gnd_net_\,
            in3 => \N__27146\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29569\,
            in2 => \_gnd_net_\,
            in3 => \N__27143\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28522\,
            in2 => \_gnd_net_\,
            in3 => \N__27251\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31093\,
            in2 => \_gnd_net_\,
            in3 => \N__27248\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28546\,
            in2 => \_gnd_net_\,
            in3 => \N__27245\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31042\,
            in2 => \_gnd_net_\,
            in3 => \N__27242\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28498\,
            in2 => \_gnd_net_\,
            in3 => \N__27239\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28900\,
            in2 => \_gnd_net_\,
            in3 => \N__27236\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27665\,
            in2 => \_gnd_net_\,
            in3 => \N__27233\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27590\,
            in2 => \_gnd_net_\,
            in3 => \N__27230\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__31428\,
            in1 => \N__27227\,
            in2 => \_gnd_net_\,
            in3 => \N__27185\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__28573\,
            in1 => \N__31422\,
            in2 => \N__27575\,
            in3 => \N__27518\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__31426\,
            in1 => \N__31043\,
            in2 => \N__31684\,
            in3 => \N__27503\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__31424\,
            in1 => \N__27491\,
            in2 => \N__29517\,
            in3 => \N__31094\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__28523\,
            in1 => \N__31795\,
            in2 => \N__27479\,
            in3 => \N__31423\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__31427\,
            in1 => \N__27457\,
            in2 => \N__28499\,
            in3 => \N__27419\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__31121\,
            in1 => \N__31421\,
            in2 => \N__27407\,
            in3 => \N__27359\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__31425\,
            in1 => \N__28547\,
            in2 => \N__31856\,
            in3 => \N__27344\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__29972\,
            in1 => \N__31511\,
            in2 => \N__27293\,
            in3 => \N__27332\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111001111"
        )
    port map (
            in0 => \N__28295\,
            in1 => \N__28157\,
            in2 => \N__27884\,
            in3 => \N__27311\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48384\,
            ce => 'H',
            sr => \N__47800\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111110"
        )
    port map (
            in0 => \N__28153\,
            in1 => \N__28296\,
            in2 => \N__27880\,
            in3 => \N__28403\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48384\,
            ce => 'H',
            sr => \N__47800\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__28293\,
            in1 => \N__28155\,
            in2 => \N__27882\,
            in3 => \N__28358\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48384\,
            ce => 'H',
            sr => \N__47800\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111110"
        )
    port map (
            in0 => \N__28154\,
            in1 => \N__28297\,
            in2 => \N__27881\,
            in3 => \N__28310\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48384\,
            ce => 'H',
            sr => \N__47800\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011111110"
        )
    port map (
            in0 => \N__28294\,
            in1 => \N__28156\,
            in2 => \N__27883\,
            in3 => \N__27782\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48384\,
            ce => 'H',
            sr => \N__47800\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__31506\,
            in1 => \N__28901\,
            in2 => \N__27731\,
            in3 => \N__27680\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27664\,
            in2 => \_gnd_net_\,
            in3 => \N__31504\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__31507\,
            in1 => \N__27650\,
            in2 => \N__27608\,
            in3 => \N__27605\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__27589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31505\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110101111101"
        )
    port map (
            in0 => \N__31508\,
            in1 => \N__28742\,
            in2 => \N__28733\,
            in3 => \N__28730\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31509\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31510\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48378\,
            ce => 'H',
            sr => \N__47804\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28569\,
            in2 => \_gnd_net_\,
            in3 => \N__31497\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31500\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28545\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29568\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31498\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31499\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28515\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__28491\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31501\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__31503\,
            in1 => \N__31070\,
            in2 => \N__28472\,
            in3 => \N__28424\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__36606\,
            in1 => \N__36471\,
            in2 => \_gnd_net_\,
            in3 => \N__36323\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31502\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28899\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30702\,
            in2 => \_gnd_net_\,
            in3 => \N__30677\,
            lcout => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__36208\,
            in1 => \N__36148\,
            in2 => \_gnd_net_\,
            in3 => \N__36122\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48363\,
            ce => \N__28843\,
            sr => \N__47821\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__32935\,
            in1 => \N__33957\,
            in2 => \_gnd_net_\,
            in3 => \N__34270\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48363\,
            ce => \N__28843\,
            sr => \N__47821\
        );

    \delay_measurement_inst.delay_hc_reg_20_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__33090\,
            in1 => \N__33499\,
            in2 => \N__30509\,
            in3 => \N__33325\,
            lcout => measured_delay_hc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48357\,
            ce => 'H',
            sr => \N__47828\
        );

    \delay_measurement_inst.delay_hc_reg_0_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__33324\,
            in1 => \N__32565\,
            in2 => \N__33522\,
            in3 => \N__33089\,
            lcout => measured_delay_hc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48357\,
            ce => 'H',
            sr => \N__47828\
        );

    \phase_controller_inst2.state_3_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__35789\,
            in1 => \N__28793\,
            in2 => \N__35822\,
            in3 => \N__33769\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48357\,
            ce => 'H',
            sr => \N__47828\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_9_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33619\,
            in1 => \N__28763\,
            in2 => \_gnd_net_\,
            in3 => \N__33321\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.N_33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_9_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110101"
        )
    port map (
            in0 => \N__33513\,
            in1 => \_gnd_net_\,
            in2 => \N__29069\,
            in3 => \N__33076\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48351\,
            ce => 'H',
            sr => \N__47837\
        );

    \delay_measurement_inst.delay_hc_reg_14_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__33512\,
            in1 => \N__29066\,
            in2 => \_gnd_net_\,
            in3 => \N__33075\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48351\,
            ce => 'H',
            sr => \N__47837\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_2_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33313\,
            in1 => \N__34039\,
            in2 => \_gnd_net_\,
            in3 => \N__29057\,
            lcout => \delay_measurement_inst.N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46379_20_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__29039\,
            in1 => \N__29017\,
            in2 => \N__29003\,
            in3 => \N__28991\,
            lcout => \delay_measurement_inst.delay_hc_reg3lt31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_18_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30748\,
            in1 => \N__28982\,
            in2 => \_gnd_net_\,
            in3 => \N__33312\,
            lcout => \delay_measurement_inst.N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__29305\,
            in1 => \N__29278\,
            in2 => \_gnd_net_\,
            in3 => \N__29226\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_303_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_24_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__33475\,
            in1 => \N__33308\,
            in2 => \N__29189\,
            in3 => \N__33042\,
            lcout => measured_delay_hc_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48342\,
            ce => 'H',
            sr => \N__47853\
        );

    \delay_measurement_inst.delay_hc_reg_4_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__33045\,
            in1 => \N__33478\,
            in2 => \_gnd_net_\,
            in3 => \N__28910\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48342\,
            ce => 'H',
            sr => \N__47853\
        );

    \delay_measurement_inst.delay_hc_reg_29_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__33477\,
            in1 => \N__30629\,
            in2 => \_gnd_net_\,
            in3 => \N__33044\,
            lcout => measured_delay_hc_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48342\,
            ce => 'H',
            sr => \N__47853\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__29309\,
            in1 => \N__29282\,
            in2 => \_gnd_net_\,
            in3 => \N__29227\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48342\,
            ce => 'H',
            sr => \N__47853\
        );

    \delay_measurement_inst.delay_hc_reg_23_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__33474\,
            in1 => \N__33307\,
            in2 => \N__29156\,
            in3 => \N__33041\,
            lcout => measured_delay_hc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48342\,
            ce => 'H',
            sr => \N__47853\
        );

    \delay_measurement_inst.delay_hc_reg_26_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__33043\,
            in1 => \N__29170\,
            in2 => \N__33326\,
            in3 => \N__33476\,
            lcout => measured_delay_hc_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48342\,
            ce => 'H',
            sr => \N__47853\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29203\,
            in1 => \N__29185\,
            in2 => \N__29174\,
            in3 => \N__29152\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__29141\,
            in1 => \N__29092\,
            in2 => \N__29123\,
            in3 => \N__30611\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_30_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30599\,
            in1 => \N__29120\,
            in2 => \_gnd_net_\,
            in3 => \N__33320\,
            lcout => \delay_measurement_inst.N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_27_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__33511\,
            in1 => \N__29102\,
            in2 => \_gnd_net_\,
            in3 => \N__33123\,
            lcout => measured_delay_hc_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48336\,
            ce => 'H',
            sr => \N__47866\
        );

    \delay_measurement_inst.delay_hc_reg_1_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__33510\,
            in1 => \N__29081\,
            in2 => \_gnd_net_\,
            in3 => \N__33122\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48336\,
            ce => 'H',
            sr => \N__47866\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42606\,
            in2 => \_gnd_net_\,
            in3 => \N__42582\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_304_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__29363\,
            in1 => \N__29345\,
            in2 => \N__47926\,
            in3 => \N__29326\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR1_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29384\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR2_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29372\,
            lcout => delay_tr_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.prev_tr_sig_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29365\,
            lcout => \delay_measurement_inst.prev_tr_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48445\,
            ce => 'H',
            sr => \N__47746\
        );

    \delay_measurement_inst.start_timer_tr_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__29364\,
            in1 => \N__29344\,
            in2 => \_gnd_net_\,
            in3 => \N__29325\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48445\,
            ce => 'H',
            sr => \N__47746\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__42634\,
            in1 => \N__42616\,
            in2 => \_gnd_net_\,
            in3 => \N__42581\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48436\,
            ce => 'H',
            sr => \N__47752\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47918\,
            in2 => \_gnd_net_\,
            in3 => \N__39277\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__30938\,
            in1 => \N__40692\,
            in2 => \_gnd_net_\,
            in3 => \N__39250\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48428\,
            ce => \N__30868\,
            sr => \N__47757\
        );

    \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111000000000"
        )
    port map (
            in0 => \N__39249\,
            in1 => \N__30937\,
            in2 => \N__40702\,
            in3 => \N__45649\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48428\,
            ce => \N__30868\,
            sr => \N__47757\
        );

    \delay_measurement_inst.delay_tr_reg_esr_2_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__40701\,
            in1 => \N__45599\,
            in2 => \N__39260\,
            in3 => \N__30936\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48418\,
            ce => \N__30870\,
            sr => \N__47766\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__29412\,
            in1 => \N__41409\,
            in2 => \_gnd_net_\,
            in3 => \N__41008\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48418\,
            ce => \N__30870\,
            sr => \N__47766\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101110"
        )
    port map (
            in0 => \N__41129\,
            in1 => \N__29413\,
            in2 => \N__41427\,
            in3 => \N__29420\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48418\,
            ce => \N__30870\,
            sr => \N__47766\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__41406\,
            in1 => \N__29409\,
            in2 => \_gnd_net_\,
            in3 => \N__41078\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48418\,
            ce => \N__30870\,
            sr => \N__47766\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__41261\,
            in1 => \N__41410\,
            in2 => \_gnd_net_\,
            in3 => \N__37257\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48418\,
            ce => \N__30870\,
            sr => \N__47766\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__41407\,
            in1 => \N__29410\,
            in2 => \_gnd_net_\,
            in3 => \N__41054\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48418\,
            ce => \N__30870\,
            sr => \N__47766\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__29411\,
            in1 => \N__41408\,
            in2 => \_gnd_net_\,
            in3 => \N__41033\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48418\,
            ce => \N__30870\,
            sr => \N__47766\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41032\,
            in1 => \N__41053\,
            in2 => \N__41009\,
            in3 => \N__41074\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10\,
            ltout => \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__41149\,
            in1 => \N__40630\,
            in2 => \N__29390\,
            in3 => \N__37245\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7\,
            ltout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29387\,
            in3 => \N__40924\,
            lcout => \delay_measurement_inst.N_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29518\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__40975\,
            in1 => \N__41111\,
            in2 => \N__40934\,
            in3 => \N__40690\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__37576\,
            in1 => \N__37511\,
            in2 => \_gnd_net_\,
            in3 => \N__37783\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38549\,
            in2 => \_gnd_net_\,
            in3 => \N__38488\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48402\,
            ce => \N__42683\,
            sr => \N__47776\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38067\,
            in2 => \_gnd_net_\,
            in3 => \N__39332\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48402\,
            ce => \N__42683\,
            sr => \N__47776\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29971\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30042\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29814\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29733\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31181\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31431\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29650\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35972\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29629\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31429\,
            in2 => \_gnd_net_\,
            in3 => \N__29608\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29850\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29760\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__31432\,
            in1 => \N__29576\,
            in2 => \N__31745\,
            in3 => \N__29546\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36014\,
            in1 => \N__29528\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30200\,
            in3 => \N__29915\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__48392\,
            ce => 'H',
            sr => \N__47785\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29912\,
            in2 => \_gnd_net_\,
            in3 => \N__29888\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__48392\,
            ce => 'H',
            sr => \N__47785\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30305\,
            in2 => \_gnd_net_\,
            in3 => \N__29864\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__48392\,
            ce => 'H',
            sr => \N__47785\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32255\,
            in2 => \_gnd_net_\,
            in3 => \N__29834\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__48392\,
            ce => 'H',
            sr => \N__47785\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29831\,
            in2 => \_gnd_net_\,
            in3 => \N__29789\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__48392\,
            ce => 'H',
            sr => \N__47785\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29786\,
            in2 => \_gnd_net_\,
            in3 => \N__29744\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__48392\,
            ce => 'H',
            sr => \N__47785\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32267\,
            in2 => \_gnd_net_\,
            in3 => \N__29711\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__48392\,
            ce => 'H',
            sr => \N__47785\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29708\,
            in2 => \_gnd_net_\,
            in3 => \N__29669\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_8\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__48388\,
            ce => 'H',
            sr => \N__47789\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30254\,
            in2 => \_gnd_net_\,
            in3 => \N__30053\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__48388\,
            ce => 'H',
            sr => \N__47789\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36770\,
            in2 => \_gnd_net_\,
            in3 => \N__30050\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__48388\,
            ce => 'H',
            sr => \N__47789\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30173\,
            in2 => \_gnd_net_\,
            in3 => \N__30020\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__48388\,
            ce => 'H',
            sr => \N__47789\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36650\,
            in2 => \_gnd_net_\,
            in3 => \N__30017\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48388\,
            ce => 'H',
            sr => \N__47789\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30006\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48388\,
            ce => 'H',
            sr => \N__47789\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36477\,
            in1 => \N__36324\,
            in2 => \N__36629\,
            in3 => \N__30101\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48388\,
            ce => 'H',
            sr => \N__47789\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29970\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \N__47792\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__36464\,
            in1 => \N__36619\,
            in2 => \N__30089\,
            in3 => \N__36328\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \N__47792\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36325\,
            in1 => \N__36468\,
            in2 => \N__36626\,
            in3 => \N__30074\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \N__47792\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__36465\,
            in1 => \N__36620\,
            in2 => \N__30065\,
            in3 => \N__36329\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \N__47792\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36326\,
            in1 => \N__36469\,
            in2 => \N__36627\,
            in3 => \N__30161\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \N__47792\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__36466\,
            in1 => \N__36621\,
            in2 => \N__30152\,
            in3 => \N__36330\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \N__47792\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36327\,
            in1 => \N__36470\,
            in2 => \N__36628\,
            in3 => \N__30140\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \N__47792\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__36467\,
            in1 => \N__36622\,
            in2 => \N__30131\,
            in3 => \N__36331\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \N__47792\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35705\,
            in2 => \N__35690\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32105\,
            in2 => \_gnd_net_\,
            in3 => \N__30092\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36026\,
            in2 => \N__32084\,
            in3 => \N__30077\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32063\,
            in2 => \_gnd_net_\,
            in3 => \N__30068\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32045\,
            in2 => \_gnd_net_\,
            in3 => \N__30056\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32012\,
            in2 => \_gnd_net_\,
            in3 => \N__30155\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31994\,
            in2 => \_gnd_net_\,
            in3 => \N__30143\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31976\,
            in2 => \_gnd_net_\,
            in3 => \N__30134\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31940\,
            in2 => \_gnd_net_\,
            in3 => \N__30119\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35651\,
            in2 => \_gnd_net_\,
            in3 => \N__30116\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35723\,
            in2 => \_gnd_net_\,
            in3 => \N__30113\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32236\,
            in2 => \_gnd_net_\,
            in3 => \N__30110\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32215\,
            in2 => \_gnd_net_\,
            in3 => \N__30107\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32194\,
            in2 => \_gnd_net_\,
            in3 => \N__30104\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32521\,
            in2 => \_gnd_net_\,
            in3 => \N__30188\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32501\,
            in2 => \_gnd_net_\,
            in3 => \N__30185\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32483\,
            in2 => \_gnd_net_\,
            in3 => \N__30182\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32465\,
            in2 => \_gnd_net_\,
            in3 => \N__30179\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32447\,
            in2 => \_gnd_net_\,
            in3 => \N__30176\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36646\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__34129\,
            in1 => \N__33922\,
            in2 => \N__30361\,
            in3 => \N__34291\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48361\,
            ce => \N__36076\,
            sr => \N__47809\
        );

    \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__34289\,
            in1 => \N__30447\,
            in2 => \N__33961\,
            in3 => \N__34128\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48361\,
            ce => \N__36076\,
            sr => \N__47809\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__34130\,
            in1 => \N__33923\,
            in2 => \N__33644\,
            in3 => \N__34292\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48361\,
            ce => \N__36076\,
            sr => \N__47809\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__30242\,
            in1 => \N__33921\,
            in2 => \_gnd_net_\,
            in3 => \N__34290\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48361\,
            ce => \N__36076\,
            sr => \N__47809\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__34288\,
            in1 => \N__30766\,
            in2 => \_gnd_net_\,
            in3 => \N__33936\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48361\,
            ce => \N__36076\,
            sr => \N__47809\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34428\,
            in1 => \N__30353\,
            in2 => \N__32936\,
            in3 => \N__34507\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto6_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__32364\,
            in1 => \N__32430\,
            in2 => \N__30451\,
            in3 => \N__30515\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35951\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30505\,
            in1 => \N__32969\,
            in2 => \N__30392\,
            in3 => \N__30295\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36668\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32674\,
            in1 => \N__30231\,
            in2 => \N__30764\,
            in3 => \N__32725\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35987\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001100"
        )
    port map (
            in0 => \N__34044\,
            in1 => \N__30398\,
            in2 => \N__32789\,
            in3 => \N__32871\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33533\,
            in1 => \N__30533\,
            in2 => \N__30527\,
            in3 => \N__30524\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34043\,
            in1 => \N__32558\,
            in2 => \N__32788\,
            in3 => \N__32870\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__30504\,
            in1 => \N__32968\,
            in2 => \N__30387\,
            in3 => \N__36123\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_5_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32357\,
            in1 => \N__30488\,
            in2 => \_gnd_net_\,
            in3 => \N__33322\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.N_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_5_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33521\,
            in2 => \N__30455\,
            in3 => \N__33059\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48345\,
            ce => 'H',
            sr => \N__47829\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__30434\,
            in1 => \N__32356\,
            in2 => \_gnd_net_\,
            in3 => \N__32425\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_21_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__33323\,
            in1 => \N__33520\,
            in2 => \N__30391\,
            in3 => \N__33058\,
            lcout => measured_delay_hc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48345\,
            ce => 'H',
            sr => \N__47829\
        );

    \delay_measurement_inst.delay_hc_reg_31_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__33516\,
            in1 => \N__33314\,
            in2 => \N__36205\,
            in3 => \N__33046\,
            lcout => measured_delay_hc_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48341\,
            ce => 'H',
            sr => \N__47838\
        );

    \delay_measurement_inst.delay_hc_reg_18_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__33047\,
            in1 => \N__33517\,
            in2 => \_gnd_net_\,
            in3 => \N__30776\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48341\,
            ce => 'H',
            sr => \N__47838\
        );

    \delay_measurement_inst.delay_hc_reg_2_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__33048\,
            in1 => \N__33518\,
            in2 => \_gnd_net_\,
            in3 => \N__30719\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48341\,
            ce => 'H',
            sr => \N__47838\
        );

    \phase_controller_inst1.state_1_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__43442\,
            in1 => \N__30713\,
            in2 => \N__43367\,
            in3 => \N__30686\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48341\,
            ce => 'H',
            sr => \N__47838\
        );

    \delay_measurement_inst.delay_hc_reg_3_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__33049\,
            in1 => \N__33519\,
            in2 => \_gnd_net_\,
            in3 => \N__30659\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48341\,
            ce => 'H',
            sr => \N__47838\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_29_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30623\,
            in1 => \N__30647\,
            in2 => \_gnd_net_\,
            in3 => \N__33318\,
            lcout => \delay_measurement_inst.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30598\,
            in2 => \_gnd_net_\,
            in3 => \N__30622\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_30_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__30605\,
            in1 => \N__33473\,
            in2 => \_gnd_net_\,
            in3 => \N__33127\,
            lcout => measured_delay_hc_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48335\,
            ce => 'H',
            sr => \N__47854\
        );

    \SB_DFF_inst_DELAY_HC1_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30587\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_13_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30575\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30821\,
            in1 => \N__30791\,
            in2 => \N__30809\,
            in3 => \N__30800\,
            lcout => \phase_controller_inst1.stoper_tr.N_248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38241\,
            in1 => \N__38686\,
            in2 => \N__38471\,
            in3 => \N__34864\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35064\,
            in2 => \_gnd_net_\,
            in3 => \N__35037\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011101"
        )
    port map (
            in0 => \N__38453\,
            in1 => \N__38545\,
            in2 => \N__30794\,
            in3 => \N__38687\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__40834\,
            in1 => \N__40935\,
            in2 => \N__41428\,
            in3 => \N__37273\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48447\,
            ce => \N__30871\,
            sr => \N__47747\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__34971\,
            in1 => \N__35169\,
            in2 => \_gnd_net_\,
            in3 => \N__35133\,
            lcout => \phase_controller_inst1.stoper_tr.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__39205\,
            in1 => \N__39327\,
            in2 => \_gnd_net_\,
            in3 => \N__34998\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38462\,
            in2 => \N__30782\,
            in3 => \N__35038\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34860\,
            in2 => \N__30779\,
            in3 => \N__38046\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48439\,
            ce => \N__42701\,
            sr => \N__47753\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__38285\,
            in1 => \N__38045\,
            in2 => \N__35113\,
            in3 => \N__34938\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48439\,
            ce => \N__42701\,
            sr => \N__47753\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010001"
        )
    port map (
            in0 => \N__40928\,
            in1 => \N__40983\,
            in2 => \N__30889\,
            in3 => \N__41121\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_ess_3_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__30933\,
            in1 => \N__40700\,
            in2 => \N__39259\,
            in3 => \N__40775\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48430\,
            ce => \N__30872\,
            sr => \N__47758\
        );

    \delay_measurement_inst.delay_tr_reg_esr_5_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__40696\,
            in1 => \N__39252\,
            in2 => \N__40727\,
            in3 => \N__30935\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48430\,
            ce => \N__30872\,
            sr => \N__47758\
        );

    \delay_measurement_inst.delay_tr_reg_esr_4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__40748\,
            in1 => \N__39251\,
            in2 => \N__40703\,
            in3 => \N__30934\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48430\,
            ce => \N__30872\,
            sr => \N__47758\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38117\,
            in1 => \N__38129\,
            in2 => \N__41456\,
            in3 => \N__30839\,
            lcout => \delay_measurement_inst.N_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__41112\,
            in1 => \N__40691\,
            in2 => \N__45650\,
            in3 => \N__40771\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__40976\,
            in1 => \N__45594\,
            in2 => \N__30842\,
            in3 => \N__40793\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41471\,
            in2 => \_gnd_net_\,
            in3 => \N__41486\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__30833\,
            in1 => \N__40847\,
            in2 => \N__41405\,
            in3 => \N__30827\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__30927\,
            in1 => \N__40833\,
            in2 => \N__30902\,
            in3 => \N__30899\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38706\,
            in1 => \N__35085\,
            in2 => \N__38583\,
            in3 => \N__38359\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38611\,
            in2 => \_gnd_net_\,
            in3 => \N__35092\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48410\,
            ce => \N__42700\,
            sr => \N__47771\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38612\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38713\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48410\,
            ce => \N__42700\,
            sr => \N__47771\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__38551\,
            in1 => \N__38472\,
            in2 => \_gnd_net_\,
            in3 => \N__38688\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111010101111"
        )
    port map (
            in0 => \N__35065\,
            in1 => \N__38497\,
            in2 => \N__30893\,
            in3 => \N__35033\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48410\,
            ce => \N__42700\,
            sr => \N__47771\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_1_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010110001000"
        )
    port map (
            in0 => \N__36376\,
            in1 => \N__36608\,
            in2 => \N__36872\,
            in3 => \N__36332\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48403\,
            ce => \N__35920\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_0_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__37440\,
            in1 => \N__37730\,
            in2 => \N__37665\,
            in3 => \N__38176\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48403\,
            ce => \N__35920\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_1_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__38177\,
            in1 => \N__37618\,
            in2 => \N__37784\,
            in3 => \N__37441\,
            lcout => \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48403\,
            ce => \N__35920\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__31400\,
            in1 => \N__31293\,
            in2 => \N__31268\,
            in3 => \N__31226\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31204\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31395\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__31401\,
            in1 => \N__31190\,
            in2 => \N__31145\,
            in3 => \N__31142\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31116\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31396\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31086\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31397\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31062\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31035\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31399\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31640\,
            in1 => \N__31013\,
            in2 => \N__31001\,
            in3 => \N__30986\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31682\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31917\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEC8M_18_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31847\,
            in1 => \N__31784\,
            in2 => \N__31744\,
            in3 => \N__31683\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31392\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__31394\,
            in1 => \N__31615\,
            in2 => \N__31571\,
            in3 => \N__31568\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__31539\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31391\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31393\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31294\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32537\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31274\,
            in2 => \N__32831\,
            in3 => \N__35679\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32090\,
            in2 => \N__33818\,
            in3 => \N__32101\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32069\,
            in2 => \N__32744\,
            in3 => \N__32080\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32062\,
            in1 => \N__32051\,
            in2 => \N__32381\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32044\,
            in1 => \N__32033\,
            in2 => \N__32327\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32000\,
            in2 => \N__32027\,
            in3 => \N__32011\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31993\,
            in1 => \N__31982\,
            in2 => \N__32693\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31961\,
            in2 => \N__32621\,
            in3 => \N__31972\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31925\,
            in2 => \N__31955\,
            in3 => \N__31936\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32180\,
            in2 => \N__32594\,
            in3 => \N__35644\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32174\,
            in2 => \N__32609\,
            in3 => \N__35719\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32237\,
            in1 => \N__32168\,
            in2 => \N__32312\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32162\,
            in2 => \N__34442\,
            in3 => \N__32216\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32141\,
            in2 => \N__32156\,
            in3 => \N__32195\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32135\,
            in2 => \N__34379\,
            in3 => \N__32522\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32129\,
            in2 => \N__32888\,
            in3 => \N__32500\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32111\,
            in2 => \N__32123\,
            in3 => \N__32482\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32282\,
            in2 => \N__32297\,
            in3 => \N__32464\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32276\,
            in2 => \N__36089\,
            in3 => \N__32446\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32270\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36704\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35936\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_1_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35826\,
            in2 => \_gnd_net_\,
            in3 => \N__35781\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36472\,
            in1 => \N__36319\,
            in2 => \N__36601\,
            in3 => \N__32243\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48373\,
            ce => 'H',
            sr => \N__47801\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36315\,
            in1 => \N__36551\,
            in2 => \N__36478\,
            in3 => \N__32222\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48373\,
            ce => 'H',
            sr => \N__47801\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36473\,
            in1 => \N__36320\,
            in2 => \N__36602\,
            in3 => \N__32201\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48373\,
            ce => 'H',
            sr => \N__47801\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36316\,
            in1 => \N__36552\,
            in2 => \N__36479\,
            in3 => \N__32528\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48373\,
            ce => 'H',
            sr => \N__47801\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36474\,
            in1 => \N__36321\,
            in2 => \N__36603\,
            in3 => \N__32507\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48373\,
            ce => 'H',
            sr => \N__47801\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100010001100"
        )
    port map (
            in0 => \N__36317\,
            in1 => \N__32489\,
            in2 => \N__36481\,
            in3 => \N__36566\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48373\,
            ce => 'H',
            sr => \N__47801\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__36475\,
            in1 => \N__32471\,
            in2 => \N__36604\,
            in3 => \N__36322\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48373\,
            ce => 'H',
            sr => \N__47801\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36318\,
            in1 => \N__36553\,
            in2 => \N__36480\,
            in3 => \N__32453\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48373\,
            ce => 'H',
            sr => \N__47801\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34294\,
            in1 => \N__32435\,
            in2 => \N__33959\,
            in3 => \N__34166\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48368\,
            ce => \N__36075\,
            sr => \N__47805\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34167\,
            in1 => \N__32365\,
            in2 => \N__34337\,
            in3 => \N__33910\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48368\,
            ce => \N__36075\,
            sr => \N__47805\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34293\,
            in1 => \N__33755\,
            in2 => \N__33958\,
            in3 => \N__34165\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48368\,
            ce => \N__36075\,
            sr => \N__47805\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__32934\,
            in1 => \N__33908\,
            in2 => \_gnd_net_\,
            in3 => \N__34296\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48368\,
            ce => \N__36075\,
            sr => \N__47805\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__33907\,
            in1 => \N__32876\,
            in2 => \_gnd_net_\,
            in3 => \N__32816\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48368\,
            ce => \N__36075\,
            sr => \N__47805\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__32817\,
            in1 => \N__33909\,
            in2 => \_gnd_net_\,
            in3 => \N__32794\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48368\,
            ce => \N__36075\,
            sr => \N__47805\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34295\,
            in1 => \N__32732\,
            in2 => \N__33960\,
            in3 => \N__34168\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48368\,
            ce => \N__36075\,
            sr => \N__47805\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34169\,
            in1 => \N__32678\,
            in2 => \N__34338\,
            in3 => \N__33911\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48368\,
            ce => \N__36075\,
            sr => \N__47805\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34172\,
            in1 => \N__33704\,
            in2 => \N__33962\,
            in3 => \N__34268\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48364\,
            ce => \N__36077\,
            sr => \N__47810\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34265\,
            in1 => \N__33927\,
            in2 => \N__33593\,
            in3 => \N__34171\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48364\,
            ce => \N__36077\,
            sr => \N__47810\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__36147\,
            in1 => \N__32579\,
            in2 => \N__36207\,
            in3 => \N__36130\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_0_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__34264\,
            in1 => \N__34170\,
            in2 => \N__32573\,
            in3 => \N__32570\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48364\,
            ce => \N__36077\,
            sr => \N__47810\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34266\,
            in1 => \N__33928\,
            in2 => \N__34508\,
            in3 => \N__34173\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48364\,
            ce => \N__36077\,
            sr => \N__47810\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34174\,
            in1 => \N__34430\,
            in2 => \N__33963\,
            in3 => \N__34269\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48364\,
            ce => \N__36077\,
            sr => \N__47810\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__34267\,
            in1 => \N__34175\,
            in2 => \N__34054\,
            in3 => \N__33935\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48364\,
            ce => \N__36077\,
            sr => \N__47810\
        );

    \phase_controller_inst1.state_3_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__33803\,
            in1 => \N__43856\,
            in2 => \N__34611\,
            in3 => \N__33773\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48358\,
            ce => 'H',
            sr => \N__47815\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33751\,
            in1 => \N__33702\,
            in2 => \N__33642\,
            in3 => \N__33574\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_22_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__33515\,
            in1 => \N__33319\,
            in2 => \N__32967\,
            in3 => \N__33128\,
            lcout => measured_delay_hc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48343\,
            ce => 'H',
            sr => \N__47839\
        );

    \current_shift_inst.timer_s1.running_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__36983\,
            in1 => \N__37004\,
            in2 => \_gnd_net_\,
            in3 => \N__34547\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48332\,
            ce => 'H',
            sr => \N__47867\
        );

    \phase_controller_inst1.S1_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34610\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48332\,
            ce => 'H',
            sr => \N__47867\
        );

    \current_shift_inst.start_timer_s1_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__34608\,
            in1 => \N__34560\,
            in2 => \_gnd_net_\,
            in3 => \N__34545\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48332\,
            ce => 'H',
            sr => \N__47867\
        );

    \current_shift_inst.stop_timer_s1_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__34546\,
            in1 => \N__34609\,
            in2 => \N__34567\,
            in3 => \N__36982\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48332\,
            ce => 'H',
            sr => \N__47867\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__37001\,
            in1 => \N__36980\,
            in2 => \_gnd_net_\,
            in3 => \N__34544\,
            lcout => \current_shift_inst.timer_s1.N_181_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43380\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48329\,
            ce => 'H',
            sr => \N__47876\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__37786\,
            in1 => \N__37677\,
            in2 => \N__37529\,
            in3 => \N__37151\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48471\,
            ce => 'H',
            sr => \N__47735\
        );

    \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_14_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37518\,
            in2 => \_gnd_net_\,
            in3 => \N__37785\,
            lcout => \phase_controller_inst2.stoper_tr.time_passed11\,
            ltout => \phase_controller_inst2.stoper_tr.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34511\,
            in3 => \N__38181\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__37792\,
            in1 => \N__37683\,
            in2 => \N__37355\,
            in3 => \N__37491\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48467\,
            ce => 'H',
            sr => \N__47738\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__37791\,
            in1 => \N__37682\,
            in2 => \N__37016\,
            in3 => \N__37490\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48467\,
            ce => 'H',
            sr => \N__47738\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__37790\,
            in1 => \N__37681\,
            in2 => \N__37097\,
            in3 => \N__37489\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48467\,
            ce => 'H',
            sr => \N__47738\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37488\,
            in1 => \N__37793\,
            in2 => \N__37685\,
            in3 => \N__36935\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48467\,
            ce => 'H',
            sr => \N__47738\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__37788\,
            in1 => \N__37527\,
            in2 => \N__37672\,
            in3 => \N__37301\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__47740\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__37524\,
            in1 => \N__37630\,
            in2 => \N__37812\,
            in3 => \N__37067\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__47740\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__37789\,
            in1 => \N__37528\,
            in2 => \N__37673\,
            in3 => \N__37127\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__47740\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__37787\,
            in1 => \N__37526\,
            in2 => \N__37671\,
            in3 => \N__37043\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__47740\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__37525\,
            in1 => \N__37631\,
            in2 => \N__37813\,
            in3 => \N__37325\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__47740\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38749\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48448\,
            ce => \N__42705\,
            sr => \N__47748\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__38275\,
            in1 => \N__38101\,
            in2 => \_gnd_net_\,
            in3 => \N__35008\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48448\,
            ce => \N__42705\,
            sr => \N__47748\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39206\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48448\,
            ce => \N__42705\,
            sr => \N__47748\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__38276\,
            in1 => \N__34978\,
            in2 => \N__38105\,
            in3 => \N__34939\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48448\,
            ce => \N__42705\,
            sr => \N__47748\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__38099\,
            in1 => \N__38274\,
            in2 => \N__35170\,
            in3 => \N__35140\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48448\,
            ce => \N__42705\,
            sr => \N__47748\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34730\,
            in2 => \N__34724\,
            in3 => \N__37830\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34703\,
            in2 => \N__34715\,
            in3 => \N__37957\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34685\,
            in2 => \N__34697\,
            in3 => \N__37930\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34679\,
            in2 => \N__38222\,
            in3 => \N__36950\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34673\,
            in2 => \N__34667\,
            in3 => \N__37906\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34643\,
            in2 => \N__34658\,
            in3 => \N__37876\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37180\,
            in1 => \N__34622\,
            in2 => \N__34637\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34829\,
            in2 => \N__34841\,
            in3 => \N__37169\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34811\,
            in2 => \N__34823\,
            in3 => \N__37142\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37852\,
            in1 => \N__34805\,
            in2 => \N__38348\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34790\,
            in2 => \N__34799\,
            in3 => \N__37381\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34769\,
            in2 => \N__34784\,
            in3 => \N__37112\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34763\,
            in2 => \N__38339\,
            in3 => \N__37082\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34757\,
            in2 => \N__38327\,
            in3 => \N__37058\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34736\,
            in2 => \N__34751\,
            in3 => \N__37034\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34922\,
            in2 => \N__42728\,
            in3 => \N__37370\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34916\,
            in2 => \N__34883\,
            in3 => \N__37343\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34910\,
            in2 => \N__34874\,
            in3 => \N__37316\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34892\,
            in2 => \N__34904\,
            in3 => \N__37214\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34886\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39127\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48421\,
            ce => \N__42709\,
            sr => \N__47767\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39079\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48421\,
            ce => \N__42709\,
            sr => \N__47767\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__38312\,
            in1 => \N__38096\,
            in2 => \_gnd_net_\,
            in3 => \N__38249\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48411\,
            ce => \N__39037\,
            sr => \N__47772\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__38094\,
            in1 => \N__34865\,
            in2 => \_gnd_net_\,
            in3 => \N__38313\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48411\,
            ce => \N__39037\,
            sr => \N__47772\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__38311\,
            in1 => \N__38095\,
            in2 => \N__35177\,
            in3 => \N__35144\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48411\,
            ce => \N__39037\,
            sr => \N__47772\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__38314\,
            in1 => \N__38097\,
            in2 => \N__35120\,
            in3 => \N__34951\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48411\,
            ce => \N__39037\,
            sr => \N__47772\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38093\,
            in2 => \_gnd_net_\,
            in3 => \N__39331\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => \N__39036\,
            sr => \N__47777\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38626\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38375\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => \N__39036\,
            sr => \N__47777\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38627\,
            in2 => \_gnd_net_\,
            in3 => \N__35096\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => \N__39036\,
            sr => \N__47777\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111010101111"
        )
    port map (
            in0 => \N__35069\,
            in1 => \N__38499\,
            in2 => \N__38641\,
            in3 => \N__35039\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => \N__39036\,
            sr => \N__47777\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__35009\,
            in1 => \N__38092\,
            in2 => \_gnd_net_\,
            in3 => \N__38307\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => \N__39036\,
            sr => \N__47777\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42764\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => \N__39036\,
            sr => \N__47777\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__38091\,
            in1 => \N__34982\,
            in2 => \N__38315\,
            in3 => \N__34952\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => \N__39036\,
            sr => \N__47777\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43562\,
            in1 => \N__43818\,
            in2 => \N__43717\,
            in3 => \N__41975\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48397\,
            ce => 'H',
            sr => \N__47779\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__43914\,
            in1 => \N__41329\,
            in2 => \_gnd_net_\,
            in3 => \N__43882\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__43565\,
            in1 => \N__43696\,
            in2 => \N__35180\,
            in3 => \N__43821\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48397\,
            ce => 'H',
            sr => \N__47779\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43815\,
            in1 => \N__43687\,
            in2 => \N__43575\,
            in3 => \N__41942\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48397\,
            ce => 'H',
            sr => \N__47779\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43563\,
            in1 => \N__43819\,
            in2 => \N__43718\,
            in3 => \N__41909\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48397\,
            ce => 'H',
            sr => \N__47779\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43816\,
            in1 => \N__43691\,
            in2 => \N__43576\,
            in3 => \N__41876\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48397\,
            ce => 'H',
            sr => \N__47779\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43564\,
            in1 => \N__43820\,
            in2 => \N__43719\,
            in3 => \N__41843\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48397\,
            ce => 'H',
            sr => \N__47779\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43817\,
            in1 => \N__43695\,
            in2 => \N__43577\,
            in3 => \N__41810\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48397\,
            ce => 'H',
            sr => \N__47779\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43776\,
            in1 => \N__43630\,
            in2 => \N__43554\,
            in3 => \N__41600\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48393\,
            ce => 'H',
            sr => \N__47786\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43517\,
            in1 => \N__43778\,
            in2 => \N__43660\,
            in3 => \N__41561\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48393\,
            ce => 'H',
            sr => \N__47786\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43777\,
            in1 => \N__43634\,
            in2 => \N__43555\,
            in3 => \N__41531\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48393\,
            ce => 'H',
            sr => \N__47786\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43629\,
            in1 => \N__43506\,
            in2 => \_gnd_net_\,
            in3 => \N__43775\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__36916\,
            in1 => \N__35683\,
            in2 => \_gnd_net_\,
            in3 => \N__36861\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__36579\,
            in1 => \N__36446\,
            in2 => \N__35693\,
            in3 => \N__36288\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48393\,
            ce => 'H',
            sr => \N__47786\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36463\,
            in1 => \N__36287\,
            in2 => \N__36609\,
            in3 => \N__35663\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48393\,
            ce => 'H',
            sr => \N__47786\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__35214\,
            in1 => \N__35355\,
            in2 => \N__35585\,
            in3 => \N__35632\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48389\,
            ce => \N__35900\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__35633\,
            in1 => \N__35574\,
            in2 => \N__35375\,
            in3 => \N__35215\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48389\,
            ce => \N__35900\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__43518\,
            in1 => \N__43804\,
            in2 => \N__43724\,
            in3 => \N__43880\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48389\,
            ce => \N__35900\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__43881\,
            in1 => \N__43716\,
            in2 => \N__43823\,
            in3 => \N__43519\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48389\,
            ce => \N__35900\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43915\,
            in2 => \_gnd_net_\,
            in3 => \N__43878\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43879\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43916\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_0_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__36459\,
            in1 => \N__36289\,
            in2 => \N__36605\,
            in3 => \N__36860\,
            lcout => \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48389\,
            ce => \N__35900\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35745\,
            in2 => \_gnd_net_\,
            in3 => \N__36807\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.start_timer_hc_RNO_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__35843\,
            in1 => \N__36550\,
            in2 => \N__35834\,
            in3 => \N__45481\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48385\,
            ce => 'H',
            sr => \N__47793\
        );

    \phase_controller_inst2.state_2_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__36808\,
            in1 => \N__35827\,
            in2 => \N__35752\,
            in3 => \N__35785\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48385\,
            ce => 'H',
            sr => \N__47793\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36549\,
            in1 => \N__36254\,
            in2 => \N__36482\,
            in3 => \N__35732\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48385\,
            ce => 'H',
            sr => \N__47793\
        );

    \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36427\,
            in2 => \_gnd_net_\,
            in3 => \N__36253\,
            lcout => \phase_controller_inst2.stoper_hc.time_passed11\,
            ltout => \phase_controller_inst2.stoper_hc.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35708\,
            in3 => \N__36849\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__36212\,
            in1 => \N__36155\,
            in2 => \_gnd_net_\,
            in3 => \N__36131\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48379\,
            ce => \N__36062\,
            sr => \N__47797\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36785\,
            in1 => \_gnd_net_\,
            in2 => \N__45966\,
            in3 => \N__45434\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45907\,
            in2 => \N__36029\,
            in3 => \N__42064\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36903\,
            in2 => \_gnd_net_\,
            in3 => \N__36850\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_0_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39167\,
            in2 => \N__39161\,
            in3 => \N__39160\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__48374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39146\,
            in2 => \_gnd_net_\,
            in3 => \N__35975\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__48374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39140\,
            in2 => \_gnd_net_\,
            in3 => \N__35954\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__48374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39407\,
            in2 => \_gnd_net_\,
            in3 => \N__35939\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__48374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39401\,
            in2 => \_gnd_net_\,
            in3 => \N__36743\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__48374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39395\,
            in2 => \_gnd_net_\,
            in3 => \N__36728\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__48374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39389\,
            in2 => \_gnd_net_\,
            in3 => \N__36707\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__48374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39359\,
            in2 => \_gnd_net_\,
            in3 => \N__36692\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__48374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36758\,
            in2 => \_gnd_net_\,
            in3 => \N__36671\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__48369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39353\,
            in2 => \_gnd_net_\,
            in3 => \N__36659\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__48369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39344\,
            in3 => \N__36656\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__48369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39662\,
            in2 => \_gnd_net_\,
            in3 => \N__36653\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__36607\,
            in1 => \N__36476\,
            in2 => \_gnd_net_\,
            in3 => \N__36296\,
            lcout => \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__49581\,
            in1 => \N__36752\,
            in2 => \_gnd_net_\,
            in3 => \N__48512\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36776\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__46462\,
            in1 => \N__42224\,
            in2 => \_gnd_net_\,
            in3 => \N__39521\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49566\,
            in1 => \N__47137\,
            in2 => \N__49280\,
            in3 => \N__47102\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48722\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48365\,
            ce => \N__47988\,
            sr => \N__47811\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46961\,
            in1 => \N__49565\,
            in2 => \N__49281\,
            in3 => \N__46193\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101111"
        )
    port map (
            in0 => \N__46192\,
            in1 => \N__49110\,
            in2 => \N__49645\,
            in3 => \N__46962\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45325\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49561\,
            in2 => \N__36746\,
            in3 => \N__48508\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49580\,
            in1 => \N__46545\,
            in2 => \N__49394\,
            in3 => \N__46505\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49588\,
            in1 => \N__49309\,
            in2 => \N__42500\,
            in3 => \N__45020\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49579\,
            in1 => \N__46926\,
            in2 => \N__49393\,
            in3 => \N__46886\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49590\,
            in1 => \N__49311\,
            in2 => \N__46783\,
            in3 => \N__46736\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49578\,
            in1 => \N__46854\,
            in2 => \N__49395\,
            in3 => \N__46814\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__49589\,
            in1 => \N__47066\,
            in2 => \N__44957\,
            in3 => \N__49310\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49577\,
            in1 => \N__44161\,
            in2 => \N__49396\,
            in3 => \N__44465\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__49587\,
            in1 => \N__44416\,
            in2 => \N__44675\,
            in3 => \N__49308\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__36806\,
            in1 => \N__36917\,
            in2 => \N__36887\,
            in3 => \N__36868\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48347\,
            ce => 'H',
            sr => \N__47830\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48705\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48338\,
            ce => \N__47954\,
            sr => \N__47848\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37002\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36981\,
            lcout => \current_shift_inst.timer_s1.N_180_i_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36962\,
            in2 => \N__37838\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_2_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_15_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37961\,
            in2 => \_gnd_net_\,
            in3 => \N__36956\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38141\,
            in2 => \N__37937\,
            in3 => \N__36953\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_15_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36949\,
            in2 => \_gnd_net_\,
            in3 => \N__36929\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37910\,
            in2 => \_gnd_net_\,
            in3 => \N__36926\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_15_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37883\,
            in2 => \_gnd_net_\,
            in3 => \N__36923\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_15_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37184\,
            in2 => \_gnd_net_\,
            in3 => \N__36920\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_15_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37165\,
            in2 => \_gnd_net_\,
            in3 => \N__37145\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37141\,
            in2 => \_gnd_net_\,
            in3 => \N__37121\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_15_3_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37856\,
            in2 => \_gnd_net_\,
            in3 => \N__37118\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37385\,
            in2 => \_gnd_net_\,
            in3 => \N__37115\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37111\,
            in2 => \_gnd_net_\,
            in3 => \N__37085\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37081\,
            in2 => \_gnd_net_\,
            in3 => \N__37061\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37057\,
            in2 => \_gnd_net_\,
            in3 => \N__37037\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37030\,
            in2 => \_gnd_net_\,
            in3 => \N__37007\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37369\,
            in2 => \_gnd_net_\,
            in3 => \N__37346\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37339\,
            in2 => \_gnd_net_\,
            in3 => \N__37319\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_15_4_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37315\,
            in2 => \_gnd_net_\,
            in3 => \N__37295\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37210\,
            in2 => \_gnd_net_\,
            in3 => \N__37292\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111110"
        )
    port map (
            in0 => \N__40829\,
            in1 => \N__37289\,
            in2 => \N__41417\,
            in3 => \N__37274\,
            lcout => \delay_measurement_inst.N_267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__37622\,
            in1 => \N__37523\,
            in2 => \_gnd_net_\,
            in3 => \N__37814\,
            lcout => \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37512\,
            in1 => \N__37803\,
            in2 => \N__37674\,
            in3 => \N__37220\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48460\,
            ce => 'H',
            sr => \N__47741\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__37802\,
            in1 => \N__37652\,
            in2 => \N__37196\,
            in3 => \N__37517\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48460\,
            ce => 'H',
            sr => \N__47741\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__37989\,
            in1 => \N__38208\,
            in2 => \N__38009\,
            in3 => \N__38183\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48460\,
            ce => 'H',
            sr => \N__47741\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__37800\,
            in1 => \N__37650\,
            in2 => \N__37973\,
            in3 => \N__37515\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48460\,
            ce => 'H',
            sr => \N__47741\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37513\,
            in1 => \N__37804\,
            in2 => \N__37675\,
            in3 => \N__37946\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48460\,
            ce => 'H',
            sr => \N__47741\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37514\,
            in1 => \N__37805\,
            in2 => \N__37676\,
            in3 => \N__37919\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48460\,
            ce => 'H',
            sr => \N__47741\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__37801\,
            in1 => \N__37651\,
            in2 => \N__37895\,
            in3 => \N__37516\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48460\,
            ce => 'H',
            sr => \N__47741\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37492\,
            in1 => \N__37810\,
            in2 => \N__37684\,
            in3 => \N__37865\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => 'H',
            sr => \N__47749\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__38210\,
            in1 => \N__37834\,
            in2 => \_gnd_net_\,
            in3 => \N__38182\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__37666\,
            in1 => \N__37493\,
            in2 => \N__37841\,
            in3 => \N__37811\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => 'H',
            sr => \N__47749\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__37809\,
            in1 => \N__37667\,
            in2 => \N__37522\,
            in3 => \N__37394\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => 'H',
            sr => \N__47749\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38642\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48440\,
            ce => \N__42687\,
            sr => \N__47754\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38643\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38590\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48440\,
            ce => \N__42687\,
            sr => \N__47754\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__38550\,
            in1 => \N__38498\,
            in2 => \_gnd_net_\,
            in3 => \N__38692\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48440\,
            ce => \N__42687\,
            sr => \N__47754\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__38297\,
            in1 => \N__38098\,
            in2 => \_gnd_net_\,
            in3 => \N__38248\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48440\,
            ce => \N__42687\,
            sr => \N__47754\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38209\,
            in2 => \_gnd_net_\,
            in3 => \N__38172\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41510\,
            in1 => \N__41519\,
            in2 => \N__41501\,
            in3 => \N__41162\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41183\,
            in1 => \N__41192\,
            in2 => \N__41174\,
            in3 => \N__41201\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42589\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38068\,
            in2 => \_gnd_net_\,
            in3 => \N__39204\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48422\,
            ce => \N__39038\,
            sr => \N__47768\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38753\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48422\,
            ce => \N__39038\,
            sr => \N__47768\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38644\,
            in2 => \_gnd_net_\,
            in3 => \N__38717\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48422\,
            ce => \N__39038\,
            sr => \N__47768\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__38693\,
            in1 => \N__38557\,
            in2 => \_gnd_net_\,
            in3 => \N__38501\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48422\,
            ce => \N__39038\,
            sr => \N__47768\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38645\,
            in2 => \_gnd_net_\,
            in3 => \N__38591\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48422\,
            ce => \N__39038\,
            sr => \N__47768\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38558\,
            in2 => \_gnd_net_\,
            in3 => \N__38500\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48422\,
            ce => \N__39038\,
            sr => \N__47768\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38411\,
            in2 => \N__38420\,
            in3 => \N__41319\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38396\,
            in2 => \N__38405\,
            in3 => \N__41305\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38381\,
            in2 => \N__38390\,
            in3 => \N__41743\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38870\,
            in2 => \N__38882\,
            in3 => \N__41713\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38852\,
            in2 => \N__38864\,
            in3 => \N__41683\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38837\,
            in2 => \N__38846\,
            in3 => \N__41650\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38822\,
            in2 => \N__38831\,
            in3 => \N__41617\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38804\,
            in2 => \N__38816\,
            in3 => \N__41584\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38789\,
            in2 => \N__38798\,
            in3 => \N__41542\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41986\,
            in1 => \N__38774\,
            in2 => \N__38783\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38759\,
            in2 => \N__38768\,
            in3 => \N__41953\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38993\,
            in2 => \N__39005\,
            in3 => \N__41920\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38975\,
            in2 => \N__38987\,
            in3 => \N__41887\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38954\,
            in2 => \N__38969\,
            in3 => \N__41854\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38936\,
            in2 => \N__38948\,
            in3 => \N__41821\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43931\,
            in1 => \N__38921\,
            in2 => \N__38930\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38915\,
            in2 => \N__39092\,
            in3 => \N__41791\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38909\,
            in2 => \N__39047\,
            in3 => \N__42109\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38888\,
            in2 => \N__38903\,
            in3 => \N__42088\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39134\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39131\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48398\,
            ce => \N__39026\,
            sr => \N__47780\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39083\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48398\,
            ce => \N__39026\,
            sr => \N__47780\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43513\,
            in1 => \N__43797\,
            in2 => \N__43720\,
            in3 => \N__41780\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48394\,
            ce => 'H',
            sr => \N__47787\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43794\,
            in1 => \N__43700\,
            in2 => \N__43556\,
            in3 => \N__42098\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48394\,
            ce => 'H',
            sr => \N__47787\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43514\,
            in1 => \N__43798\,
            in2 => \N__43721\,
            in3 => \N__42074\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48394\,
            ce => 'H',
            sr => \N__47787\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43795\,
            in1 => \N__43704\,
            in2 => \N__43557\,
            in3 => \N__41771\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48394\,
            ce => 'H',
            sr => \N__47787\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010000010"
        )
    port map (
            in0 => \N__41726\,
            in1 => \N__43526\,
            in2 => \N__43722\,
            in3 => \N__43800\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48394\,
            ce => 'H',
            sr => \N__47787\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43796\,
            in1 => \N__43708\,
            in2 => \N__43558\,
            in3 => \N__41696\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48394\,
            ce => 'H',
            sr => \N__47787\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43515\,
            in1 => \N__43799\,
            in2 => \N__43723\,
            in3 => \N__41666\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48394\,
            ce => 'H',
            sr => \N__47787\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__41633\,
            in1 => \N__43516\,
            in2 => \N__43822\,
            in3 => \N__43712\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48394\,
            ce => 'H',
            sr => \N__47787\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46694\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45231\,
            in1 => \N__49741\,
            in2 => \N__49391\,
            in3 => \N__44794\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49744\,
            in1 => \N__44412\,
            in2 => \N__49388\,
            in3 => \N__44671\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48686\,
            in1 => \N__42492\,
            in2 => \_gnd_net_\,
            in3 => \N__45018\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__45019\,
            in1 => \N__49292\,
            in2 => \N__42499\,
            in3 => \N__49749\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49750\,
            in1 => \N__47069\,
            in2 => \N__49390\,
            in3 => \N__44956\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49743\,
            in1 => \N__44536\,
            in2 => \N__49389\,
            in3 => \N__44627\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__45232\,
            in1 => \N__49742\,
            in2 => \N__49392\,
            in3 => \N__44795\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__42236\,
            in1 => \N__39536\,
            in2 => \_gnd_net_\,
            in3 => \N__46459\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__39509\,
            in1 => \N__42212\,
            in2 => \_gnd_net_\,
            in3 => \N__46460\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__46461\,
            in1 => \N__39497\,
            in2 => \_gnd_net_\,
            in3 => \N__42200\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_7_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__39247\,
            in1 => \N__40637\,
            in2 => \N__39326\,
            in3 => \N__39286\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48386\,
            ce => 'H',
            sr => \N__47794\
        );

    \delay_measurement_inst.delay_tr_reg_8_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__39287\,
            in1 => \N__39248\,
            in2 => \N__39189\,
            in3 => \N__41153\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48386\,
            ce => 'H',
            sr => \N__47794\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__39464\,
            in1 => \N__42167\,
            in2 => \_gnd_net_\,
            in3 => \N__46438\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46439\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.N_1318_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__39452\,
            in1 => \N__42158\,
            in2 => \_gnd_net_\,
            in3 => \N__46440\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__46441\,
            in1 => \N__39620\,
            in2 => \_gnd_net_\,
            in3 => \N__42149\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__42140\,
            in1 => \N__39605\,
            in2 => \_gnd_net_\,
            in3 => \N__46442\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__46443\,
            in1 => \N__39581\,
            in2 => \_gnd_net_\,
            in3 => \N__42278\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__39566\,
            in1 => \N__42269\,
            in2 => \_gnd_net_\,
            in3 => \N__46444\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__46445\,
            in1 => \N__39551\,
            in2 => \_gnd_net_\,
            in3 => \N__42260\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39383\,
            in2 => \N__42043\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46403\,
            in2 => \N__46349\,
            in3 => \N__45396\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45397\,
            in1 => \N__39377\,
            in2 => \N__49195\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48975\,
            in2 => \N__39371\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46562\,
            in2 => \N__49196\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48979\,
            in2 => \N__42350\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39440\,
            in2 => \N__49197\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48983\,
            in2 => \N__42176\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48984\,
            in2 => \N__42305\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48994\,
            in2 => \N__42359\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39428\,
            in2 => \N__49201\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39422\,
            in2 => \N__49198\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42329\,
            in2 => \N__49202\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39413\,
            in2 => \N__49199\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42395\,
            in2 => \N__49203\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39485\,
            in2 => \N__49200\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49204\,
            in2 => \N__42407\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39479\,
            in2 => \N__49356\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49208\,
            in2 => \N__39473\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42284\,
            in2 => \N__49357\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49212\,
            in2 => \N__42455\,
            in3 => \N__39455\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49802\,
            in2 => \N__49358\,
            in3 => \N__39443\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49216\,
            in2 => \N__39629\,
            in3 => \N__39608\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42386\,
            in2 => \N__49359\,
            in3 => \N__39593\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49220\,
            in2 => \N__39590\,
            in3 => \N__39569\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42365\,
            in2 => \N__49360\,
            in3 => \N__39554\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49224\,
            in2 => \N__42425\,
            in3 => \N__39539\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42461\,
            in2 => \N__49361\,
            in3 => \N__39524\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42371\,
            in2 => \N__49428\,
            in3 => \N__39512\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42446\,
            in2 => \N__49362\,
            in3 => \N__39500\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42439\,
            in2 => \N__49429\,
            in3 => \N__39488\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_0_11_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010100110101"
        )
    port map (
            in0 => \N__42185\,
            in1 => \N__49811\,
            in2 => \N__46466\,
            in3 => \N__39665\,
            lcout => \current_shift_inst.control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39817\,
            in2 => \N__48545\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__48352\,
            ce => \N__48008\,
            sr => \N__47822\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39796\,
            in2 => \N__46393\,
            in3 => \N__39650\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__48352\,
            ce => \N__48008\,
            sr => \N__47822\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39818\,
            in2 => \N__39772\,
            in3 => \N__39647\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__48352\,
            ce => \N__48008\,
            sr => \N__47822\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39797\,
            in2 => \N__39745\,
            in3 => \N__39644\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__48352\,
            ce => \N__48008\,
            sr => \N__47822\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40039\,
            in2 => \N__39773\,
            in3 => \N__39641\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__48352\,
            ce => \N__48008\,
            sr => \N__47822\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40015\,
            in2 => \N__39746\,
            in3 => \N__39638\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__48352\,
            ce => \N__48008\,
            sr => \N__47822\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40040\,
            in2 => \N__39992\,
            in3 => \N__39635\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__48352\,
            ce => \N__48008\,
            sr => \N__47822\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40016\,
            in2 => \N__39962\,
            in3 => \N__39632\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__48352\,
            ce => \N__48008\,
            sr => \N__47822\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39991\,
            in2 => \N__39931\,
            in3 => \N__39692\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__48348\,
            ce => \N__47995\,
            sr => \N__47831\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39961\,
            in2 => \N__39901\,
            in3 => \N__39689\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__48348\,
            ce => \N__47995\,
            sr => \N__47831\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39874\,
            in2 => \N__39932\,
            in3 => \N__39686\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__48348\,
            ce => \N__47995\,
            sr => \N__47831\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39853\,
            in2 => \N__39902\,
            in3 => \N__39683\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__48348\,
            ce => \N__47995\,
            sr => \N__47831\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39875\,
            in2 => \N__40258\,
            in3 => \N__39680\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__48348\,
            ce => \N__47995\,
            sr => \N__47831\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39854\,
            in2 => \N__40231\,
            in3 => \N__39677\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__48348\,
            ce => \N__47995\,
            sr => \N__47831\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40201\,
            in2 => \N__40259\,
            in3 => \N__39674\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__48348\,
            ce => \N__47995\,
            sr => \N__47831\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40174\,
            in2 => \N__40232\,
            in3 => \N__39671\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__48348\,
            ce => \N__47995\,
            sr => \N__47831\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40202\,
            in2 => \N__40144\,
            in3 => \N__39668\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__48344\,
            ce => \N__47987\,
            sr => \N__47840\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40175\,
            in2 => \N__40114\,
            in3 => \N__39719\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__48344\,
            ce => \N__47987\,
            sr => \N__47840\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40084\,
            in2 => \N__40145\,
            in3 => \N__39716\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__48344\,
            ce => \N__47987\,
            sr => \N__47840\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40063\,
            in2 => \N__40115\,
            in3 => \N__39713\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__48344\,
            ce => \N__47987\,
            sr => \N__47840\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40085\,
            in2 => \N__40609\,
            in3 => \N__39710\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__48344\,
            ce => \N__47987\,
            sr => \N__47840\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40064\,
            in2 => \N__40579\,
            in3 => \N__39707\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__48344\,
            ce => \N__47987\,
            sr => \N__47840\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40552\,
            in2 => \N__40610\,
            in3 => \N__39704\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__48344\,
            ce => \N__47987\,
            sr => \N__47840\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40525\,
            in2 => \N__40580\,
            in3 => \N__39701\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__48344\,
            ce => \N__47987\,
            sr => \N__47840\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40553\,
            in2 => \N__40498\,
            in3 => \N__39698\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__48339\,
            ce => \N__47994\,
            sr => \N__47849\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40526\,
            in2 => \N__40468\,
            in3 => \N__39695\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__48339\,
            ce => \N__47994\,
            sr => \N__47849\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40439\,
            in2 => \N__40499\,
            in3 => \N__39833\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__48339\,
            ce => \N__47994\,
            sr => \N__47849\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40295\,
            in2 => \N__40469\,
            in3 => \N__39830\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__48339\,
            ce => \N__47994\,
            sr => \N__47849\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39827\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40380\,
            in1 => \N__48531\,
            in2 => \_gnd_net_\,
            in3 => \N__39824\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__48337\,
            ce => \N__40277\,
            sr => \N__47855\
        );

    \current_shift_inst.timer_s1.counter_1_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40375\,
            in1 => \N__46380\,
            in2 => \_gnd_net_\,
            in3 => \N__39821\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__48337\,
            ce => \N__40277\,
            sr => \N__47855\
        );

    \current_shift_inst.timer_s1.counter_2_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40381\,
            in1 => \N__39816\,
            in2 => \_gnd_net_\,
            in3 => \N__39800\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__48337\,
            ce => \N__40277\,
            sr => \N__47855\
        );

    \current_shift_inst.timer_s1.counter_3_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40376\,
            in1 => \N__39790\,
            in2 => \_gnd_net_\,
            in3 => \N__39776\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__48337\,
            ce => \N__40277\,
            sr => \N__47855\
        );

    \current_shift_inst.timer_s1.counter_4_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40382\,
            in1 => \N__39765\,
            in2 => \_gnd_net_\,
            in3 => \N__39749\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__48337\,
            ce => \N__40277\,
            sr => \N__47855\
        );

    \current_shift_inst.timer_s1.counter_5_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40377\,
            in1 => \N__39738\,
            in2 => \_gnd_net_\,
            in3 => \N__39722\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__48337\,
            ce => \N__40277\,
            sr => \N__47855\
        );

    \current_shift_inst.timer_s1.counter_6_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40379\,
            in1 => \N__40033\,
            in2 => \_gnd_net_\,
            in3 => \N__40019\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__48337\,
            ce => \N__40277\,
            sr => \N__47855\
        );

    \current_shift_inst.timer_s1.counter_7_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40378\,
            in1 => \N__40009\,
            in2 => \_gnd_net_\,
            in3 => \N__39995\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__48337\,
            ce => \N__40277\,
            sr => \N__47855\
        );

    \current_shift_inst.timer_s1.counter_8_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40386\,
            in1 => \N__39981\,
            in2 => \_gnd_net_\,
            in3 => \N__39965\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__48334\,
            ce => \N__40276\,
            sr => \N__47861\
        );

    \current_shift_inst.timer_s1.counter_9_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40412\,
            in1 => \N__39951\,
            in2 => \_gnd_net_\,
            in3 => \N__39935\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__48334\,
            ce => \N__40276\,
            sr => \N__47861\
        );

    \current_shift_inst.timer_s1.counter_10_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40383\,
            in1 => \N__39919\,
            in2 => \_gnd_net_\,
            in3 => \N__39905\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__48334\,
            ce => \N__40276\,
            sr => \N__47861\
        );

    \current_shift_inst.timer_s1.counter_11_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40409\,
            in1 => \N__39894\,
            in2 => \_gnd_net_\,
            in3 => \N__39878\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__48334\,
            ce => \N__40276\,
            sr => \N__47861\
        );

    \current_shift_inst.timer_s1.counter_12_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40384\,
            in1 => \N__39873\,
            in2 => \_gnd_net_\,
            in3 => \N__39857\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__48334\,
            ce => \N__40276\,
            sr => \N__47861\
        );

    \current_shift_inst.timer_s1.counter_13_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40410\,
            in1 => \N__39852\,
            in2 => \_gnd_net_\,
            in3 => \N__39836\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__48334\,
            ce => \N__40276\,
            sr => \N__47861\
        );

    \current_shift_inst.timer_s1.counter_14_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40385\,
            in1 => \N__40251\,
            in2 => \_gnd_net_\,
            in3 => \N__40235\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__48334\,
            ce => \N__40276\,
            sr => \N__47861\
        );

    \current_shift_inst.timer_s1.counter_15_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40411\,
            in1 => \N__40219\,
            in2 => \_gnd_net_\,
            in3 => \N__40205\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__48334\,
            ce => \N__40276\,
            sr => \N__47861\
        );

    \current_shift_inst.timer_s1.counter_16_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40401\,
            in1 => \N__40194\,
            in2 => \_gnd_net_\,
            in3 => \N__40178\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_15_27_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__48333\,
            ce => \N__40275\,
            sr => \N__47868\
        );

    \current_shift_inst.timer_s1.counter_17_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40405\,
            in1 => \N__40167\,
            in2 => \_gnd_net_\,
            in3 => \N__40148\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__48333\,
            ce => \N__40275\,
            sr => \N__47868\
        );

    \current_shift_inst.timer_s1.counter_18_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40402\,
            in1 => \N__40132\,
            in2 => \_gnd_net_\,
            in3 => \N__40118\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__48333\,
            ce => \N__40275\,
            sr => \N__47868\
        );

    \current_shift_inst.timer_s1.counter_19_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40406\,
            in1 => \N__40102\,
            in2 => \_gnd_net_\,
            in3 => \N__40088\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__48333\,
            ce => \N__40275\,
            sr => \N__47868\
        );

    \current_shift_inst.timer_s1.counter_20_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40403\,
            in1 => \N__40083\,
            in2 => \_gnd_net_\,
            in3 => \N__40067\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__48333\,
            ce => \N__40275\,
            sr => \N__47868\
        );

    \current_shift_inst.timer_s1.counter_21_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40407\,
            in1 => \N__40057\,
            in2 => \_gnd_net_\,
            in3 => \N__40043\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__48333\,
            ce => \N__40275\,
            sr => \N__47868\
        );

    \current_shift_inst.timer_s1.counter_22_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40404\,
            in1 => \N__40597\,
            in2 => \_gnd_net_\,
            in3 => \N__40583\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__48333\,
            ce => \N__40275\,
            sr => \N__47868\
        );

    \current_shift_inst.timer_s1.counter_23_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40408\,
            in1 => \N__40572\,
            in2 => \_gnd_net_\,
            in3 => \N__40556\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__48333\,
            ce => \N__40275\,
            sr => \N__47868\
        );

    \current_shift_inst.timer_s1.counter_24_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40413\,
            in1 => \N__40545\,
            in2 => \_gnd_net_\,
            in3 => \N__40529\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_15_28_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__48331\,
            ce => \N__40274\,
            sr => \N__47872\
        );

    \current_shift_inst.timer_s1.counter_25_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40417\,
            in1 => \N__40518\,
            in2 => \_gnd_net_\,
            in3 => \N__40502\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__48331\,
            ce => \N__40274\,
            sr => \N__47872\
        );

    \current_shift_inst.timer_s1.counter_26_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40414\,
            in1 => \N__40486\,
            in2 => \_gnd_net_\,
            in3 => \N__40472\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__48331\,
            ce => \N__40274\,
            sr => \N__47872\
        );

    \current_shift_inst.timer_s1.counter_27_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40418\,
            in1 => \N__40456\,
            in2 => \_gnd_net_\,
            in3 => \N__40442\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__48331\,
            ce => \N__40274\,
            sr => \N__47872\
        );

    \current_shift_inst.timer_s1.counter_28_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40415\,
            in1 => \N__40435\,
            in2 => \_gnd_net_\,
            in3 => \N__40421\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__48331\,
            ce => \N__40274\,
            sr => \N__47872\
        );

    \current_shift_inst.timer_s1.counter_29_LC_15_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__40291\,
            in1 => \N__40416\,
            in2 => \_gnd_net_\,
            in3 => \N__40298\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48331\,
            ce => \N__40274\,
            sr => \N__47872\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__41256\,
            in1 => \N__40764\,
            in2 => \N__41232\,
            in3 => \N__45595\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__41280\,
            in1 => \N__40872\,
            in2 => \N__40850\,
            in3 => \N__40786\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__41257\,
            in1 => \N__41281\,
            in2 => \N__41233\,
            in3 => \N__40873\,
            lcout => \delay_measurement_inst.N_265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40741\,
            in2 => \_gnd_net_\,
            in3 => \N__40717\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_287_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45667\,
            in2 => \N__42544\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_16_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__48450\,
            ce => \N__45564\,
            sr => \N__47750\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45616\,
            in2 => \N__42520\,
            in3 => \N__40730\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__48450\,
            ce => \N__45564\,
            sr => \N__47750\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42942\,
            in2 => \N__42545\,
            in3 => \N__40706\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__48450\,
            ce => \N__45564\,
            sr => \N__47750\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42924\,
            in2 => \N__42521\,
            in3 => \N__40640\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__48450\,
            ce => \N__45564\,
            sr => \N__47750\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42943\,
            in2 => \N__42907\,
            in3 => \N__40613\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__48450\,
            ce => \N__45564\,
            sr => \N__47750\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42925\,
            in2 => \N__42883\,
            in3 => \N__41132\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__48450\,
            ce => \N__45564\,
            sr => \N__47750\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42860\,
            in2 => \N__42908\,
            in3 => \N__41081\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__48450\,
            ce => \N__45564\,
            sr => \N__47750\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42836\,
            in2 => \N__42884\,
            in3 => \N__41057\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__48450\,
            ce => \N__45564\,
            sr => \N__47750\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42859\,
            in2 => \N__42811\,
            in3 => \N__41036\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__48441\,
            ce => \N__45565\,
            sr => \N__47755\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42835\,
            in2 => \N__42787\,
            in3 => \N__41012\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__48441\,
            ce => \N__45565\,
            sr => \N__47755\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43125\,
            in2 => \N__42812\,
            in3 => \N__40988\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__48441\,
            ce => \N__45565\,
            sr => \N__47755\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43107\,
            in2 => \N__42788\,
            in3 => \N__40940\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__48441\,
            ce => \N__45565\,
            sr => \N__47755\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43126\,
            in2 => \N__43090\,
            in3 => \N__40883\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__48441\,
            ce => \N__45565\,
            sr => \N__47755\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43108\,
            in2 => \N__43066\,
            in3 => \N__40853\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__48441\,
            ce => \N__45565\,
            sr => \N__47755\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43043\,
            in2 => \N__43091\,
            in3 => \N__41264\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__48441\,
            ce => \N__45565\,
            sr => \N__47755\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43019\,
            in2 => \N__43067\,
            in3 => \N__41237\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__48441\,
            ce => \N__45565\,
            sr => \N__47755\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43042\,
            in2 => \N__42994\,
            in3 => \N__41204\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__48431\,
            ce => \N__45567\,
            sr => \N__47759\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43018\,
            in2 => \N__42970\,
            in3 => \N__41195\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__48431\,
            ce => \N__45567\,
            sr => \N__47759\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43320\,
            in2 => \N__42995\,
            in3 => \N__41186\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__48431\,
            ce => \N__45567\,
            sr => \N__47759\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43302\,
            in2 => \N__42971\,
            in3 => \N__41177\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__48431\,
            ce => \N__45567\,
            sr => \N__47759\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43321\,
            in2 => \N__43285\,
            in3 => \N__41165\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__48431\,
            ce => \N__45567\,
            sr => \N__47759\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43303\,
            in2 => \N__43261\,
            in3 => \N__41156\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__48431\,
            ce => \N__45567\,
            sr => \N__47759\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43238\,
            in2 => \N__43286\,
            in3 => \N__41513\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__48431\,
            ce => \N__45567\,
            sr => \N__47759\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43214\,
            in2 => \N__43262\,
            in3 => \N__41504\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__48431\,
            ce => \N__45567\,
            sr => \N__47759\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43237\,
            in2 => \N__43189\,
            in3 => \N__41489\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__48423\,
            ce => \N__45569\,
            sr => \N__47769\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43213\,
            in2 => \N__43165\,
            in3 => \N__41474\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__48423\,
            ce => \N__45569\,
            sr => \N__47769\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43141\,
            in2 => \N__43190\,
            in3 => \N__41459\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__48423\,
            ce => \N__45569\,
            sr => \N__47769\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43984\,
            in2 => \N__43166\,
            in3 => \N__41441\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__48423\,
            ce => \N__45569\,
            sr => \N__47769\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41438\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48423\,
            ce => \N__45569\,
            sr => \N__47769\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41342\,
            in2 => \N__41330\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41306\,
            in2 => \_gnd_net_\,
            in3 => \N__41762\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41759\,
            in2 => \N__41747\,
            in3 => \N__41717\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41714\,
            in2 => \_gnd_net_\,
            in3 => \N__41687\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41684\,
            in2 => \_gnd_net_\,
            in3 => \N__41657\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41654\,
            in2 => \_gnd_net_\,
            in3 => \N__41624\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41621\,
            in2 => \_gnd_net_\,
            in3 => \N__41588\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41585\,
            in2 => \_gnd_net_\,
            in3 => \N__41549\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41546\,
            in2 => \_gnd_net_\,
            in3 => \N__41522\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41993\,
            in2 => \_gnd_net_\,
            in3 => \N__41963\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41960\,
            in2 => \_gnd_net_\,
            in3 => \N__41930\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41927\,
            in2 => \_gnd_net_\,
            in3 => \N__41897\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41894\,
            in2 => \_gnd_net_\,
            in3 => \N__41864\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41861\,
            in2 => \_gnd_net_\,
            in3 => \N__41831\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41828\,
            in2 => \_gnd_net_\,
            in3 => \N__41798\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43930\,
            in2 => \_gnd_net_\,
            in3 => \N__41795\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41792\,
            in2 => \_gnd_net_\,
            in3 => \N__41774\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42110\,
            in2 => \_gnd_net_\,
            in3 => \N__42092\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42089\,
            in2 => \_gnd_net_\,
            in3 => \N__42077\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42068\,
            in2 => \N__42044\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46319\,
            in2 => \N__46354\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42014\,
            in2 => \N__49349\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49170\,
            in2 => \N__44138\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44177\,
            in2 => \N__49350\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49174\,
            in2 => \N__44219\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41999\,
            in2 => \N__49351\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49178\,
            in2 => \N__44276\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49179\,
            in2 => \N__44591\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44423\,
            in2 => \N__49352\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49183\,
            in2 => \N__42131\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44486\,
            in2 => \N__49353\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49187\,
            in2 => \N__44288\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42122\,
            in2 => \N__49354\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49191\,
            in2 => \N__44129\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42116\,
            in2 => \N__49355\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49068\,
            in2 => \N__44306\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42380\,
            in2 => \N__49272\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49072\,
            in2 => \N__42317\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44582\,
            in2 => \N__49273\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49076\,
            in2 => \N__45359\,
            in3 => \N__42161\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48782\,
            in2 => \N__49274\,
            in3 => \N__42152\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49080\,
            in2 => \N__42341\,
            in3 => \N__42143\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44294\,
            in2 => \N__49275\,
            in3 => \N__42134\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42323\,
            in2 => \N__49276\,
            in3 => \N__42272\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49087\,
            in2 => \N__42296\,
            in3 => \N__42263\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42416\,
            in2 => \N__49277\,
            in3 => \N__42254\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49091\,
            in2 => \N__42251\,
            in3 => \N__42227\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47021\,
            in2 => \N__49278\,
            in3 => \N__42215\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49095\,
            in2 => \N__45341\,
            in3 => \N__42203\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42440\,
            in2 => \N__49279\,
            in3 => \N__42191\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_2_11_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__49790\,
            in1 => \N__49099\,
            in2 => \_gnd_net_\,
            in3 => \N__42188\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49618\,
            in1 => \N__44205\,
            in2 => \N__49285\,
            in3 => \N__44757\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49106\,
            in1 => \N__49620\,
            in2 => \N__44378\,
            in3 => \N__44703\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49617\,
            in1 => \N__44262\,
            in2 => \N__49284\,
            in3 => \N__44817\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49103\,
            in1 => \N__49623\,
            in2 => \N__46931\,
            in3 => \N__46882\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49621\,
            in1 => \N__47437\,
            in2 => \N__49282\,
            in3 => \N__47386\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49104\,
            in1 => \N__49624\,
            in2 => \N__46550\,
            in3 => \N__46501\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49622\,
            in1 => \N__46855\,
            in2 => \N__49283\,
            in3 => \N__46810\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49105\,
            in1 => \N__49619\,
            in2 => \N__45191\,
            in3 => \N__44737\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49249\,
            in1 => \N__49757\,
            in2 => \N__46267\,
            in3 => \N__46219\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__49754\,
            in1 => \N__46701\,
            in2 => \N__46648\,
            in3 => \N__49256\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__49250\,
            in1 => \N__47356\,
            in2 => \N__47318\,
            in3 => \N__49756\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49753\,
            in1 => \N__49254\,
            in2 => \N__44576\,
            in3 => \N__44898\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44334\,
            in1 => \N__49751\,
            in2 => \N__49378\,
            in3 => \N__44976\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47426\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49248\,
            in1 => \N__49755\,
            in2 => \N__45287\,
            in3 => \N__45114\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49752\,
            in1 => \N__49255\,
            in2 => \N__46784\,
            in3 => \N__46732\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49763\,
            in1 => \N__47008\,
            in2 => \N__49379\,
            in3 => \N__46979\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49266\,
            in1 => \N__49762\,
            in2 => \N__46268\,
            in3 => \N__46218\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44193\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47282\,
            in1 => \N__49761\,
            in2 => \N__49381\,
            in3 => \N__47255\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49765\,
            in1 => \N__47227\,
            in2 => \N__49380\,
            in3 => \N__47186\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44237\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__49764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47159\,
            lcout => \current_shift_inst.un4_control_input_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44151\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44355\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44317\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__49785\,
            in1 => \N__47317\,
            in2 => \N__49433\,
            in3 => \N__47349\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44396\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46593\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42477\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49786\,
            in1 => \N__47136\,
            in2 => \N__49432\,
            in3 => \N__47095\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46754\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48754\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44507\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46904\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46832\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46238\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46990\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47336\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44556\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46521\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47115\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42760\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48472\,
            ce => \N__42710\,
            sr => \N__47736\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__42641\,
            in1 => \N__42620\,
            in2 => \_gnd_net_\,
            in3 => \N__42590\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_305_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44113\,
            in1 => \N__45666\,
            in2 => \_gnd_net_\,
            in3 => \N__42551\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__48461\,
            ce => \N__43955\,
            sr => \N__47742\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44117\,
            in1 => \N__45615\,
            in2 => \_gnd_net_\,
            in3 => \N__42548\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__48461\,
            ce => \N__43955\,
            sr => \N__47742\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44114\,
            in1 => \N__42543\,
            in2 => \_gnd_net_\,
            in3 => \N__42524\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__48461\,
            ce => \N__43955\,
            sr => \N__47742\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44118\,
            in1 => \N__42519\,
            in2 => \_gnd_net_\,
            in3 => \N__42947\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__48461\,
            ce => \N__43955\,
            sr => \N__47742\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44115\,
            in1 => \N__42944\,
            in2 => \_gnd_net_\,
            in3 => \N__42929\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__48461\,
            ce => \N__43955\,
            sr => \N__47742\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44119\,
            in1 => \N__42926\,
            in2 => \_gnd_net_\,
            in3 => \N__42911\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__48461\,
            ce => \N__43955\,
            sr => \N__47742\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44116\,
            in1 => \N__42906\,
            in2 => \_gnd_net_\,
            in3 => \N__42887\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__48461\,
            ce => \N__43955\,
            sr => \N__47742\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44120\,
            in1 => \N__42882\,
            in2 => \_gnd_net_\,
            in3 => \N__42863\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__48461\,
            ce => \N__43955\,
            sr => \N__47742\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44057\,
            in1 => \N__42858\,
            in2 => \_gnd_net_\,
            in3 => \N__42839\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__48451\,
            ce => \N__43965\,
            sr => \N__47751\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44080\,
            in1 => \N__42834\,
            in2 => \_gnd_net_\,
            in3 => \N__42815\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__48451\,
            ce => \N__43965\,
            sr => \N__47751\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44054\,
            in1 => \N__42810\,
            in2 => \_gnd_net_\,
            in3 => \N__42791\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__48451\,
            ce => \N__43965\,
            sr => \N__47751\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44077\,
            in1 => \N__42786\,
            in2 => \_gnd_net_\,
            in3 => \N__42767\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__48451\,
            ce => \N__43965\,
            sr => \N__47751\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44055\,
            in1 => \N__43127\,
            in2 => \_gnd_net_\,
            in3 => \N__43112\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__48451\,
            ce => \N__43965\,
            sr => \N__47751\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44078\,
            in1 => \N__43109\,
            in2 => \_gnd_net_\,
            in3 => \N__43094\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__48451\,
            ce => \N__43965\,
            sr => \N__47751\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44056\,
            in1 => \N__43089\,
            in2 => \_gnd_net_\,
            in3 => \N__43070\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__48451\,
            ce => \N__43965\,
            sr => \N__47751\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44079\,
            in1 => \N__43065\,
            in2 => \_gnd_net_\,
            in3 => \N__43046\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__48451\,
            ce => \N__43965\,
            sr => \N__47751\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44091\,
            in1 => \N__43041\,
            in2 => \_gnd_net_\,
            in3 => \N__43022\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__48442\,
            ce => \N__43973\,
            sr => \N__47756\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44085\,
            in1 => \N__43017\,
            in2 => \_gnd_net_\,
            in3 => \N__42998\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__48442\,
            ce => \N__43973\,
            sr => \N__47756\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44092\,
            in1 => \N__42993\,
            in2 => \_gnd_net_\,
            in3 => \N__42974\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__48442\,
            ce => \N__43973\,
            sr => \N__47756\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44086\,
            in1 => \N__42969\,
            in2 => \_gnd_net_\,
            in3 => \N__42950\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__48442\,
            ce => \N__43973\,
            sr => \N__47756\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44093\,
            in1 => \N__43322\,
            in2 => \_gnd_net_\,
            in3 => \N__43307\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__48442\,
            ce => \N__43973\,
            sr => \N__47756\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44087\,
            in1 => \N__43304\,
            in2 => \_gnd_net_\,
            in3 => \N__43289\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__48442\,
            ce => \N__43973\,
            sr => \N__47756\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44094\,
            in1 => \N__43284\,
            in2 => \_gnd_net_\,
            in3 => \N__43265\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__48442\,
            ce => \N__43973\,
            sr => \N__47756\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44088\,
            in1 => \N__43260\,
            in2 => \_gnd_net_\,
            in3 => \N__43241\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__48442\,
            ce => \N__43973\,
            sr => \N__47756\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44081\,
            in1 => \N__43236\,
            in2 => \_gnd_net_\,
            in3 => \N__43217\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__48432\,
            ce => \N__43969\,
            sr => \N__47760\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44089\,
            in1 => \N__43212\,
            in2 => \_gnd_net_\,
            in3 => \N__43193\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__48432\,
            ce => \N__43969\,
            sr => \N__47760\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44082\,
            in1 => \N__43188\,
            in2 => \_gnd_net_\,
            in3 => \N__43169\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__48432\,
            ce => \N__43969\,
            sr => \N__47760\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44090\,
            in1 => \N__43164\,
            in2 => \_gnd_net_\,
            in3 => \N__43145\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__48432\,
            ce => \N__43969\,
            sr => \N__47760\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44083\,
            in1 => \N__43142\,
            in2 => \_gnd_net_\,
            in3 => \N__43130\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__48432\,
            ce => \N__43969\,
            sr => \N__47760\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__43985\,
            in1 => \N__44084\,
            in2 => \_gnd_net_\,
            in3 => \N__43988\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48432\,
            ce => \N__43969\,
            sr => \N__47760\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43561\,
            in1 => \N__43826\,
            in2 => \N__43683\,
            in3 => \N__43937\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48424\,
            ce => 'H',
            sr => \N__47770\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43559\,
            in2 => \_gnd_net_\,
            in3 => \N__43824\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed11\,
            ltout => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010111000"
        )
    port map (
            in0 => \N__43402\,
            in1 => \N__43448\,
            in2 => \N__43892\,
            in3 => \N__43889\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48424\,
            ce => 'H',
            sr => \N__47770\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43401\,
            in2 => \_gnd_net_\,
            in3 => \N__43333\,
            lcout => \phase_controller_inst1.state_RNI7NN7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__43825\,
            in1 => \N__43640\,
            in2 => \_gnd_net_\,
            in3 => \N__43560\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__43435\,
            in1 => \N__43403\,
            in2 => \N__43388\,
            in3 => \N__43334\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48412\,
            ce => 'H',
            sr => \N__47773\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48687\,
            in1 => \N__44263\,
            in2 => \_gnd_net_\,
            in3 => \N__44821\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__44759\,
            in1 => \N__49748\,
            in2 => \N__44210\,
            in3 => \N__49443\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49747\,
            in1 => \N__49427\,
            in2 => \N__44267\,
            in3 => \N__44822\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48670\,
            in1 => \N__46612\,
            in2 => \_gnd_net_\,
            in3 => \N__46579\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48689\,
            in1 => \N__44206\,
            in2 => \_gnd_net_\,
            in3 => \N__44758\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49746\,
            in1 => \N__46613\,
            in2 => \N__49450\,
            in3 => \N__46580\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48688\,
            in1 => \N__45236\,
            in2 => \_gnd_net_\,
            in3 => \N__44788\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48669\,
            in1 => \N__44167\,
            in2 => \_gnd_net_\,
            in3 => \N__44460\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__44461\,
            in1 => \N__49745\,
            in2 => \N__44171\,
            in3 => \N__49423\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__44978\,
            in1 => \N__49776\,
            in2 => \N__44339\,
            in3 => \N__49439\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49775\,
            in1 => \N__44377\,
            in2 => \N__49454\,
            in3 => \N__44705\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44417\,
            in1 => \N__48673\,
            in2 => \_gnd_net_\,
            in3 => \N__44664\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48672\,
            in1 => \N__44376\,
            in2 => \_gnd_net_\,
            in3 => \N__44704\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47068\,
            in1 => \N__48676\,
            in2 => \_gnd_net_\,
            in3 => \N__44943\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48675\,
            in1 => \N__44335\,
            in2 => \_gnd_net_\,
            in3 => \N__44977\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44535\,
            in1 => \N__48674\,
            in2 => \_gnd_net_\,
            in3 => \N__44622\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48671\,
            in1 => \N__45189\,
            in2 => \_gnd_net_\,
            in3 => \N__44738\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44572\,
            in1 => \N__49780\,
            in2 => \N__49457\,
            in3 => \N__44902\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49782\,
            in1 => \N__45283\,
            in2 => \N__49434\,
            in3 => \N__45116\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__47390\,
            in1 => \N__49779\,
            in2 => \N__47438\,
            in3 => \N__49401\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49777\,
            in1 => \N__45190\,
            in2 => \N__49435\,
            in3 => \N__44736\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__46649\,
            in1 => \N__49781\,
            in2 => \N__46706\,
            in3 => \N__49402\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__48665\,
            in1 => \_gnd_net_\,
            in2 => \N__44903\,
            in3 => \N__44571\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__44626\,
            in1 => \N__49778\,
            in2 => \N__44540\,
            in3 => \N__49400\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48666\,
            in1 => \N__45282\,
            in2 => \_gnd_net_\,
            in3 => \N__45115\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46361\,
            in2 => \N__45326\,
            in3 => \N__45324\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46937\,
            in2 => \_gnd_net_\,
            in3 => \N__44480\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44477\,
            in2 => \_gnd_net_\,
            in3 => \N__44441\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44438\,
            in2 => \_gnd_net_\,
            in3 => \N__44426\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44831\,
            in2 => \_gnd_net_\,
            in3 => \N__44798\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45200\,
            in2 => \_gnd_net_\,
            in3 => \N__44771\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44768\,
            in2 => \_gnd_net_\,
            in3 => \N__44741\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45149\,
            in2 => \_gnd_net_\,
            in3 => \N__44717\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44714\,
            in2 => \_gnd_net_\,
            in3 => \N__44687\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44684\,
            in2 => \_gnd_net_\,
            in3 => \N__44642\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44639\,
            in2 => \_gnd_net_\,
            in3 => \N__44603\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44600\,
            in2 => \_gnd_net_\,
            in3 => \N__44594\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45029\,
            in2 => \_gnd_net_\,
            in3 => \N__44993\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44990\,
            in2 => \_gnd_net_\,
            in3 => \N__44960\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47027\,
            in2 => \_gnd_net_\,
            in3 => \N__44918\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44915\,
            in2 => \_gnd_net_\,
            in3 => \N__44882\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44879\,
            in2 => \_gnd_net_\,
            in3 => \N__44870\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44867\,
            in2 => \_gnd_net_\,
            in3 => \N__44855\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44852\,
            in2 => \_gnd_net_\,
            in3 => \N__44837\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46475\,
            in2 => \_gnd_net_\,
            in3 => \N__44834\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45140\,
            in2 => \_gnd_net_\,
            in3 => \N__45131\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45128\,
            in2 => \_gnd_net_\,
            in3 => \N__45119\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45245\,
            in2 => \_gnd_net_\,
            in3 => \N__45098\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45095\,
            in2 => \_gnd_net_\,
            in3 => \N__45083\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45080\,
            in2 => \_gnd_net_\,
            in3 => \N__45071\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45068\,
            in2 => \_gnd_net_\,
            in3 => \N__45059\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45056\,
            in2 => \_gnd_net_\,
            in3 => \N__45044\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45041\,
            in2 => \_gnd_net_\,
            in3 => \N__45032\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45677\,
            in2 => \_gnd_net_\,
            in3 => \N__45365\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45362\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49784\,
            in1 => \N__47288\,
            in2 => \N__49431\,
            in3 => \N__47254\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49766\,
            in1 => \N__49377\,
            in2 => \N__47228\,
            in3 => \N__47185\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48495\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__48496\,
            in1 => \_gnd_net_\,
            in2 => \N__45290\,
            in3 => \N__48575\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45281\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45227\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45171\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47205\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45668\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48473\,
            ce => \N__45566\,
            sr => \N__47737\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45617\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48468\,
            ce => \N__45568\,
            sr => \N__47739\
        );

    \phase_controller_inst1.state_4_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45510\,
            in2 => \_gnd_net_\,
            in3 => \N__45458\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48433\,
            ce => 'H',
            sr => \N__47761\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45433\,
            in2 => \N__45404\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46277\,
            in2 => \N__46148\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46172\,
            in2 => \N__46116\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45377\,
            in2 => \N__46149\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45371\,
            in2 => \N__46117\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45722\,
            in2 => \N__46150\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45716\,
            in2 => \N__46118\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45710\,
            in2 => \N__46151\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46129\,
            in2 => \N__45704\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45695\,
            in2 => \N__46147\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45689\,
            in2 => \N__46113\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45683\,
            in2 => \N__46145\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47369\,
            in2 => \N__46114\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46068\,
            in2 => \N__45752\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45740\,
            in2 => \N__46115\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45734\,
            in2 => \N__46146\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45728\,
            in2 => \N__46119\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46715\,
            in2 => \N__46059\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46793\,
            in2 => \N__46120\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46622\,
            in2 => \N__46060\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47237\,
            in2 => \N__46121\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48731\,
            in2 => \N__46061\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46865\,
            in2 => \N__46122\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46094\,
            in2 => \N__46160\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46484\,
            in2 => \N__46035\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46199\,
            in2 => \N__46039\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47297\,
            in2 => \N__46036\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47078\,
            in2 => \N__46040\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49820\,
            in2 => \N__46037\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47168\,
            in2 => \N__46041\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47147\,
            in2 => \N__46038\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49783\,
            in2 => \_gnd_net_\,
            in3 => \N__46469\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__49707\,
            in1 => \N__46303\,
            in2 => \N__46355\,
            in3 => \N__46291\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46394\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48390\,
            ce => \N__48017\,
            sr => \N__47790\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46289\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__46292\,
            in1 => \N__49708\,
            in2 => \N__46307\,
            in3 => \N__46353\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__48604\,
            in1 => \N__46302\,
            in2 => \_gnd_net_\,
            in3 => \N__46290\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49709\,
            in1 => \N__46266\,
            in2 => \_gnd_net_\,
            in3 => \N__46220\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46964\,
            in1 => \N__48605\,
            in2 => \_gnd_net_\,
            in3 => \N__46183\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46963\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48668\,
            in1 => \N__46930\,
            in2 => \_gnd_net_\,
            in3 => \N__46881\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48606\,
            in1 => \N__46856\,
            in2 => \_gnd_net_\,
            in3 => \N__46809\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48667\,
            in1 => \N__46782\,
            in2 => \_gnd_net_\,
            in3 => \N__46731\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48607\,
            in1 => \N__46702\,
            in2 => \_gnd_net_\,
            in3 => \N__46638\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49710\,
            in1 => \N__46611\,
            in2 => \N__49455\,
            in3 => \N__46578\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48608\,
            in1 => \N__46546\,
            in2 => \_gnd_net_\,
            in3 => \N__46500\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47286\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48658\,
            in1 => \N__47427\,
            in2 => \_gnd_net_\,
            in3 => \N__47385\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49738\,
            in1 => \N__47357\,
            in2 => \_gnd_net_\,
            in3 => \N__47313\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__47287\,
            in1 => \_gnd_net_\,
            in2 => \N__48685\,
            in3 => \N__47253\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49739\,
            in1 => \N__47223\,
            in2 => \_gnd_net_\,
            in3 => \N__47184\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49740\,
            in2 => \_gnd_net_\,
            in3 => \N__47158\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49737\,
            in1 => \N__47138\,
            in2 => \_gnd_net_\,
            in3 => \N__47094\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47067\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__46978\,
            in1 => \N__49735\,
            in2 => \N__47009\,
            in3 => \N__49370\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49733\,
            in1 => \N__47004\,
            in2 => \_gnd_net_\,
            in3 => \N__46977\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_1_11_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49736\,
            in2 => \_gnd_net_\,
            in3 => \N__49369\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49732\,
            in1 => \N__48769\,
            in2 => \N__49430\,
            in3 => \N__48742\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__48743\,
            in1 => \N__49734\,
            in2 => \N__49456\,
            in3 => \N__48770\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48603\,
            in1 => \N__48768\,
            in2 => \_gnd_net_\,
            in3 => \N__48741\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48721\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48375\,
            ce => \N__48012\,
            sr => \N__47802\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48544\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48370\,
            ce => \N__48016\,
            sr => \N__47806\
        );
end \INTERFACE\;
