// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 13 2025 23:22:37

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    rgb_g,
    T01,
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    clock_output,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output rgb_g;
    output T01;
    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output clock_output;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__48639;
    wire N__48638;
    wire N__48637;
    wire N__48628;
    wire N__48627;
    wire N__48626;
    wire N__48619;
    wire N__48618;
    wire N__48617;
    wire N__48610;
    wire N__48609;
    wire N__48608;
    wire N__48601;
    wire N__48600;
    wire N__48599;
    wire N__48592;
    wire N__48591;
    wire N__48590;
    wire N__48583;
    wire N__48582;
    wire N__48581;
    wire N__48574;
    wire N__48573;
    wire N__48572;
    wire N__48565;
    wire N__48564;
    wire N__48563;
    wire N__48556;
    wire N__48555;
    wire N__48554;
    wire N__48547;
    wire N__48546;
    wire N__48545;
    wire N__48538;
    wire N__48537;
    wire N__48536;
    wire N__48529;
    wire N__48528;
    wire N__48527;
    wire N__48520;
    wire N__48519;
    wire N__48518;
    wire N__48511;
    wire N__48510;
    wire N__48509;
    wire N__48502;
    wire N__48501;
    wire N__48500;
    wire N__48493;
    wire N__48492;
    wire N__48491;
    wire N__48484;
    wire N__48483;
    wire N__48482;
    wire N__48465;
    wire N__48464;
    wire N__48463;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48449;
    wire N__48448;
    wire N__48445;
    wire N__48442;
    wire N__48439;
    wire N__48436;
    wire N__48431;
    wire N__48426;
    wire N__48425;
    wire N__48422;
    wire N__48421;
    wire N__48418;
    wire N__48415;
    wire N__48412;
    wire N__48405;
    wire N__48402;
    wire N__48401;
    wire N__48400;
    wire N__48397;
    wire N__48394;
    wire N__48391;
    wire N__48388;
    wire N__48385;
    wire N__48378;
    wire N__48377;
    wire N__48376;
    wire N__48373;
    wire N__48370;
    wire N__48367;
    wire N__48362;
    wire N__48359;
    wire N__48358;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48342;
    wire N__48341;
    wire N__48340;
    wire N__48339;
    wire N__48338;
    wire N__48337;
    wire N__48336;
    wire N__48335;
    wire N__48334;
    wire N__48333;
    wire N__48332;
    wire N__48331;
    wire N__48330;
    wire N__48329;
    wire N__48328;
    wire N__48327;
    wire N__48326;
    wire N__48325;
    wire N__48324;
    wire N__48323;
    wire N__48322;
    wire N__48315;
    wire N__48314;
    wire N__48311;
    wire N__48310;
    wire N__48309;
    wire N__48308;
    wire N__48307;
    wire N__48306;
    wire N__48305;
    wire N__48302;
    wire N__48301;
    wire N__48300;
    wire N__48299;
    wire N__48298;
    wire N__48297;
    wire N__48296;
    wire N__48295;
    wire N__48294;
    wire N__48293;
    wire N__48292;
    wire N__48291;
    wire N__48290;
    wire N__48289;
    wire N__48288;
    wire N__48287;
    wire N__48286;
    wire N__48285;
    wire N__48284;
    wire N__48279;
    wire N__48272;
    wire N__48269;
    wire N__48268;
    wire N__48267;
    wire N__48266;
    wire N__48265;
    wire N__48264;
    wire N__48263;
    wire N__48262;
    wire N__48261;
    wire N__48260;
    wire N__48259;
    wire N__48258;
    wire N__48257;
    wire N__48256;
    wire N__48255;
    wire N__48254;
    wire N__48253;
    wire N__48252;
    wire N__48251;
    wire N__48250;
    wire N__48249;
    wire N__48248;
    wire N__48247;
    wire N__48234;
    wire N__48231;
    wire N__48230;
    wire N__48229;
    wire N__48228;
    wire N__48227;
    wire N__48226;
    wire N__48225;
    wire N__48220;
    wire N__48217;
    wire N__48214;
    wire N__48201;
    wire N__48196;
    wire N__48193;
    wire N__48192;
    wire N__48191;
    wire N__48190;
    wire N__48189;
    wire N__48188;
    wire N__48187;
    wire N__48186;
    wire N__48185;
    wire N__48184;
    wire N__48173;
    wire N__48166;
    wire N__48163;
    wire N__48152;
    wire N__48143;
    wire N__48138;
    wire N__48135;
    wire N__48132;
    wire N__48121;
    wire N__48120;
    wire N__48119;
    wire N__48118;
    wire N__48115;
    wire N__48106;
    wire N__48101;
    wire N__48092;
    wire N__48081;
    wire N__48078;
    wire N__48075;
    wire N__48074;
    wire N__48073;
    wire N__48060;
    wire N__48057;
    wire N__48050;
    wire N__48045;
    wire N__48044;
    wire N__48043;
    wire N__48042;
    wire N__48041;
    wire N__48034;
    wire N__48031;
    wire N__48026;
    wire N__48019;
    wire N__48014;
    wire N__48011;
    wire N__48004;
    wire N__47999;
    wire N__47996;
    wire N__47993;
    wire N__47988;
    wire N__47985;
    wire N__47978;
    wire N__47971;
    wire N__47966;
    wire N__47957;
    wire N__47954;
    wire N__47947;
    wire N__47944;
    wire N__47939;
    wire N__47928;
    wire N__47925;
    wire N__47914;
    wire N__47895;
    wire N__47892;
    wire N__47891;
    wire N__47886;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47876;
    wire N__47875;
    wire N__47874;
    wire N__47873;
    wire N__47870;
    wire N__47869;
    wire N__47866;
    wire N__47863;
    wire N__47862;
    wire N__47861;
    wire N__47858;
    wire N__47855;
    wire N__47852;
    wire N__47851;
    wire N__47850;
    wire N__47849;
    wire N__47848;
    wire N__47847;
    wire N__47844;
    wire N__47843;
    wire N__47842;
    wire N__47841;
    wire N__47840;
    wire N__47839;
    wire N__47838;
    wire N__47837;
    wire N__47836;
    wire N__47835;
    wire N__47834;
    wire N__47833;
    wire N__47832;
    wire N__47831;
    wire N__47830;
    wire N__47829;
    wire N__47828;
    wire N__47827;
    wire N__47826;
    wire N__47825;
    wire N__47824;
    wire N__47823;
    wire N__47822;
    wire N__47821;
    wire N__47820;
    wire N__47819;
    wire N__47816;
    wire N__47815;
    wire N__47812;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47802;
    wire N__47799;
    wire N__47796;
    wire N__47793;
    wire N__47784;
    wire N__47781;
    wire N__47780;
    wire N__47779;
    wire N__47778;
    wire N__47777;
    wire N__47770;
    wire N__47761;
    wire N__47752;
    wire N__47743;
    wire N__47736;
    wire N__47735;
    wire N__47732;
    wire N__47729;
    wire N__47726;
    wire N__47717;
    wire N__47714;
    wire N__47711;
    wire N__47708;
    wire N__47705;
    wire N__47702;
    wire N__47699;
    wire N__47696;
    wire N__47685;
    wire N__47676;
    wire N__47671;
    wire N__47664;
    wire N__47661;
    wire N__47656;
    wire N__47653;
    wire N__47648;
    wire N__47645;
    wire N__47640;
    wire N__47635;
    wire N__47632;
    wire N__47623;
    wire N__47618;
    wire N__47613;
    wire N__47610;
    wire N__47607;
    wire N__47604;
    wire N__47601;
    wire N__47598;
    wire N__47583;
    wire N__47580;
    wire N__47577;
    wire N__47576;
    wire N__47573;
    wire N__47570;
    wire N__47567;
    wire N__47564;
    wire N__47559;
    wire N__47556;
    wire N__47555;
    wire N__47554;
    wire N__47553;
    wire N__47552;
    wire N__47551;
    wire N__47550;
    wire N__47549;
    wire N__47548;
    wire N__47547;
    wire N__47546;
    wire N__47545;
    wire N__47544;
    wire N__47543;
    wire N__47542;
    wire N__47541;
    wire N__47540;
    wire N__47539;
    wire N__47538;
    wire N__47537;
    wire N__47536;
    wire N__47535;
    wire N__47534;
    wire N__47533;
    wire N__47532;
    wire N__47531;
    wire N__47530;
    wire N__47529;
    wire N__47528;
    wire N__47527;
    wire N__47526;
    wire N__47525;
    wire N__47524;
    wire N__47523;
    wire N__47522;
    wire N__47521;
    wire N__47520;
    wire N__47519;
    wire N__47518;
    wire N__47517;
    wire N__47516;
    wire N__47515;
    wire N__47514;
    wire N__47513;
    wire N__47512;
    wire N__47511;
    wire N__47510;
    wire N__47509;
    wire N__47508;
    wire N__47507;
    wire N__47506;
    wire N__47505;
    wire N__47504;
    wire N__47503;
    wire N__47502;
    wire N__47501;
    wire N__47500;
    wire N__47499;
    wire N__47498;
    wire N__47497;
    wire N__47496;
    wire N__47495;
    wire N__47494;
    wire N__47493;
    wire N__47492;
    wire N__47491;
    wire N__47490;
    wire N__47489;
    wire N__47488;
    wire N__47487;
    wire N__47486;
    wire N__47485;
    wire N__47484;
    wire N__47483;
    wire N__47482;
    wire N__47481;
    wire N__47480;
    wire N__47479;
    wire N__47478;
    wire N__47477;
    wire N__47476;
    wire N__47475;
    wire N__47474;
    wire N__47473;
    wire N__47472;
    wire N__47471;
    wire N__47470;
    wire N__47469;
    wire N__47468;
    wire N__47467;
    wire N__47466;
    wire N__47465;
    wire N__47464;
    wire N__47463;
    wire N__47462;
    wire N__47461;
    wire N__47460;
    wire N__47459;
    wire N__47458;
    wire N__47457;
    wire N__47456;
    wire N__47455;
    wire N__47454;
    wire N__47453;
    wire N__47452;
    wire N__47451;
    wire N__47450;
    wire N__47449;
    wire N__47448;
    wire N__47447;
    wire N__47446;
    wire N__47445;
    wire N__47444;
    wire N__47443;
    wire N__47442;
    wire N__47441;
    wire N__47440;
    wire N__47439;
    wire N__47438;
    wire N__47437;
    wire N__47436;
    wire N__47435;
    wire N__47434;
    wire N__47433;
    wire N__47432;
    wire N__47431;
    wire N__47430;
    wire N__47429;
    wire N__47428;
    wire N__47427;
    wire N__47426;
    wire N__47425;
    wire N__47424;
    wire N__47423;
    wire N__47422;
    wire N__47421;
    wire N__47420;
    wire N__47419;
    wire N__47418;
    wire N__47417;
    wire N__47416;
    wire N__47413;
    wire N__47412;
    wire N__47127;
    wire N__47124;
    wire N__47123;
    wire N__47122;
    wire N__47121;
    wire N__47118;
    wire N__47115;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47103;
    wire N__47100;
    wire N__47099;
    wire N__47098;
    wire N__47095;
    wire N__47094;
    wire N__47093;
    wire N__47092;
    wire N__47091;
    wire N__47090;
    wire N__47089;
    wire N__47088;
    wire N__47087;
    wire N__47086;
    wire N__47085;
    wire N__47084;
    wire N__47083;
    wire N__47082;
    wire N__47081;
    wire N__47080;
    wire N__47079;
    wire N__47078;
    wire N__47077;
    wire N__47076;
    wire N__47075;
    wire N__47074;
    wire N__47073;
    wire N__47072;
    wire N__47071;
    wire N__47070;
    wire N__47069;
    wire N__47068;
    wire N__47067;
    wire N__47066;
    wire N__47065;
    wire N__47064;
    wire N__47063;
    wire N__47062;
    wire N__47061;
    wire N__47060;
    wire N__47059;
    wire N__47058;
    wire N__47057;
    wire N__47056;
    wire N__47055;
    wire N__47054;
    wire N__47053;
    wire N__47052;
    wire N__47051;
    wire N__47050;
    wire N__47049;
    wire N__47048;
    wire N__47047;
    wire N__47046;
    wire N__47045;
    wire N__47044;
    wire N__47043;
    wire N__47042;
    wire N__47041;
    wire N__47040;
    wire N__47039;
    wire N__47038;
    wire N__47037;
    wire N__47036;
    wire N__47035;
    wire N__47034;
    wire N__47033;
    wire N__47032;
    wire N__47031;
    wire N__47030;
    wire N__47029;
    wire N__47028;
    wire N__47027;
    wire N__47026;
    wire N__47025;
    wire N__47024;
    wire N__47023;
    wire N__47022;
    wire N__47021;
    wire N__47020;
    wire N__47019;
    wire N__47018;
    wire N__47017;
    wire N__47016;
    wire N__47015;
    wire N__47014;
    wire N__47013;
    wire N__47012;
    wire N__47011;
    wire N__47010;
    wire N__47009;
    wire N__47008;
    wire N__47007;
    wire N__47006;
    wire N__47005;
    wire N__47004;
    wire N__47003;
    wire N__47002;
    wire N__47001;
    wire N__47000;
    wire N__46999;
    wire N__46998;
    wire N__46997;
    wire N__46996;
    wire N__46995;
    wire N__46994;
    wire N__46993;
    wire N__46992;
    wire N__46991;
    wire N__46990;
    wire N__46989;
    wire N__46988;
    wire N__46987;
    wire N__46986;
    wire N__46985;
    wire N__46984;
    wire N__46983;
    wire N__46982;
    wire N__46981;
    wire N__46980;
    wire N__46979;
    wire N__46978;
    wire N__46977;
    wire N__46976;
    wire N__46975;
    wire N__46974;
    wire N__46973;
    wire N__46972;
    wire N__46971;
    wire N__46970;
    wire N__46969;
    wire N__46968;
    wire N__46967;
    wire N__46966;
    wire N__46965;
    wire N__46964;
    wire N__46963;
    wire N__46962;
    wire N__46961;
    wire N__46960;
    wire N__46959;
    wire N__46958;
    wire N__46957;
    wire N__46956;
    wire N__46955;
    wire N__46662;
    wire N__46659;
    wire N__46656;
    wire N__46655;
    wire N__46652;
    wire N__46651;
    wire N__46650;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46626;
    wire N__46623;
    wire N__46620;
    wire N__46613;
    wire N__46608;
    wire N__46605;
    wire N__46604;
    wire N__46601;
    wire N__46598;
    wire N__46593;
    wire N__46592;
    wire N__46589;
    wire N__46588;
    wire N__46587;
    wire N__46584;
    wire N__46581;
    wire N__46578;
    wire N__46573;
    wire N__46568;
    wire N__46563;
    wire N__46560;
    wire N__46559;
    wire N__46558;
    wire N__46555;
    wire N__46550;
    wire N__46547;
    wire N__46546;
    wire N__46543;
    wire N__46540;
    wire N__46537;
    wire N__46536;
    wire N__46533;
    wire N__46530;
    wire N__46527;
    wire N__46524;
    wire N__46521;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46502;
    wire N__46501;
    wire N__46498;
    wire N__46493;
    wire N__46488;
    wire N__46487;
    wire N__46484;
    wire N__46481;
    wire N__46476;
    wire N__46475;
    wire N__46470;
    wire N__46467;
    wire N__46466;
    wire N__46463;
    wire N__46460;
    wire N__46457;
    wire N__46456;
    wire N__46455;
    wire N__46452;
    wire N__46449;
    wire N__46446;
    wire N__46443;
    wire N__46440;
    wire N__46435;
    wire N__46434;
    wire N__46433;
    wire N__46430;
    wire N__46425;
    wire N__46420;
    wire N__46413;
    wire N__46410;
    wire N__46407;
    wire N__46404;
    wire N__46401;
    wire N__46398;
    wire N__46395;
    wire N__46392;
    wire N__46389;
    wire N__46388;
    wire N__46385;
    wire N__46382;
    wire N__46377;
    wire N__46374;
    wire N__46373;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46357;
    wire N__46354;
    wire N__46353;
    wire N__46350;
    wire N__46345;
    wire N__46342;
    wire N__46335;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46319;
    wire N__46318;
    wire N__46315;
    wire N__46312;
    wire N__46309;
    wire N__46304;
    wire N__46301;
    wire N__46300;
    wire N__46295;
    wire N__46292;
    wire N__46287;
    wire N__46284;
    wire N__46281;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46271;
    wire N__46268;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46248;
    wire N__46245;
    wire N__46240;
    wire N__46237;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46217;
    wire N__46214;
    wire N__46211;
    wire N__46210;
    wire N__46205;
    wire N__46204;
    wire N__46201;
    wire N__46198;
    wire N__46195;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46176;
    wire N__46173;
    wire N__46172;
    wire N__46171;
    wire N__46168;
    wire N__46165;
    wire N__46162;
    wire N__46157;
    wire N__46152;
    wire N__46149;
    wire N__46148;
    wire N__46147;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46117;
    wire N__46114;
    wire N__46107;
    wire N__46104;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46082;
    wire N__46081;
    wire N__46080;
    wire N__46079;
    wire N__46078;
    wire N__46077;
    wire N__46076;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46044;
    wire N__46043;
    wire N__46038;
    wire N__46037;
    wire N__46034;
    wire N__46031;
    wire N__46028;
    wire N__46023;
    wire N__46022;
    wire N__46019;
    wire N__46014;
    wire N__46013;
    wire N__46010;
    wire N__46007;
    wire N__46004;
    wire N__45999;
    wire N__45998;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45984;
    wire N__45981;
    wire N__45978;
    wire N__45977;
    wire N__45974;
    wire N__45971;
    wire N__45968;
    wire N__45963;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45953;
    wire N__45950;
    wire N__45949;
    wire N__45946;
    wire N__45943;
    wire N__45940;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45926;
    wire N__45925;
    wire N__45922;
    wire N__45919;
    wire N__45916;
    wire N__45913;
    wire N__45906;
    wire N__45905;
    wire N__45902;
    wire N__45899;
    wire N__45894;
    wire N__45891;
    wire N__45888;
    wire N__45885;
    wire N__45882;
    wire N__45879;
    wire N__45876;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45863;
    wire N__45860;
    wire N__45855;
    wire N__45854;
    wire N__45851;
    wire N__45848;
    wire N__45845;
    wire N__45840;
    wire N__45839;
    wire N__45836;
    wire N__45835;
    wire N__45832;
    wire N__45827;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45800;
    wire N__45797;
    wire N__45794;
    wire N__45789;
    wire N__45786;
    wire N__45783;
    wire N__45782;
    wire N__45781;
    wire N__45778;
    wire N__45773;
    wire N__45768;
    wire N__45767;
    wire N__45764;
    wire N__45761;
    wire N__45758;
    wire N__45755;
    wire N__45750;
    wire N__45749;
    wire N__45744;
    wire N__45741;
    wire N__45738;
    wire N__45737;
    wire N__45734;
    wire N__45731;
    wire N__45726;
    wire N__45725;
    wire N__45720;
    wire N__45717;
    wire N__45716;
    wire N__45711;
    wire N__45708;
    wire N__45707;
    wire N__45702;
    wire N__45699;
    wire N__45696;
    wire N__45693;
    wire N__45692;
    wire N__45687;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45677;
    wire N__45672;
    wire N__45669;
    wire N__45666;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45654;
    wire N__45651;
    wire N__45650;
    wire N__45649;
    wire N__45648;
    wire N__45645;
    wire N__45640;
    wire N__45637;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45617;
    wire N__45612;
    wire N__45611;
    wire N__45608;
    wire N__45605;
    wire N__45600;
    wire N__45597;
    wire N__45596;
    wire N__45595;
    wire N__45592;
    wire N__45587;
    wire N__45586;
    wire N__45581;
    wire N__45578;
    wire N__45575;
    wire N__45572;
    wire N__45569;
    wire N__45566;
    wire N__45561;
    wire N__45558;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45546;
    wire N__45543;
    wire N__45542;
    wire N__45541;
    wire N__45538;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45521;
    wire N__45520;
    wire N__45517;
    wire N__45514;
    wire N__45511;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45495;
    wire N__45494;
    wire N__45493;
    wire N__45490;
    wire N__45485;
    wire N__45480;
    wire N__45479;
    wire N__45478;
    wire N__45475;
    wire N__45472;
    wire N__45467;
    wire N__45462;
    wire N__45461;
    wire N__45456;
    wire N__45453;
    wire N__45450;
    wire N__45447;
    wire N__45444;
    wire N__45441;
    wire N__45438;
    wire N__45435;
    wire N__45432;
    wire N__45429;
    wire N__45428;
    wire N__45427;
    wire N__45424;
    wire N__45421;
    wire N__45416;
    wire N__45411;
    wire N__45410;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45398;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45384;
    wire N__45381;
    wire N__45378;
    wire N__45377;
    wire N__45374;
    wire N__45371;
    wire N__45370;
    wire N__45369;
    wire N__45364;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45350;
    wire N__45345;
    wire N__45344;
    wire N__45341;
    wire N__45340;
    wire N__45337;
    wire N__45334;
    wire N__45331;
    wire N__45326;
    wire N__45323;
    wire N__45318;
    wire N__45317;
    wire N__45316;
    wire N__45313;
    wire N__45310;
    wire N__45307;
    wire N__45302;
    wire N__45301;
    wire N__45298;
    wire N__45295;
    wire N__45292;
    wire N__45289;
    wire N__45284;
    wire N__45279;
    wire N__45276;
    wire N__45275;
    wire N__45272;
    wire N__45271;
    wire N__45268;
    wire N__45265;
    wire N__45262;
    wire N__45255;
    wire N__45252;
    wire N__45249;
    wire N__45246;
    wire N__45243;
    wire N__45242;
    wire N__45241;
    wire N__45238;
    wire N__45233;
    wire N__45228;
    wire N__45227;
    wire N__45224;
    wire N__45223;
    wire N__45220;
    wire N__45215;
    wire N__45210;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45194;
    wire N__45193;
    wire N__45188;
    wire N__45185;
    wire N__45182;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45172;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45158;
    wire N__45155;
    wire N__45152;
    wire N__45147;
    wire N__45146;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45134;
    wire N__45133;
    wire N__45132;
    wire N__45129;
    wire N__45122;
    wire N__45117;
    wire N__45116;
    wire N__45113;
    wire N__45110;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45096;
    wire N__45093;
    wire N__45092;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45080;
    wire N__45079;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45065;
    wire N__45060;
    wire N__45057;
    wire N__45056;
    wire N__45053;
    wire N__45052;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45040;
    wire N__45037;
    wire N__45032;
    wire N__45027;
    wire N__45024;
    wire N__45021;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45011;
    wire N__45010;
    wire N__45007;
    wire N__45004;
    wire N__45001;
    wire N__44996;
    wire N__44991;
    wire N__44990;
    wire N__44987;
    wire N__44984;
    wire N__44983;
    wire N__44980;
    wire N__44977;
    wire N__44976;
    wire N__44973;
    wire N__44968;
    wire N__44965;
    wire N__44962;
    wire N__44957;
    wire N__44952;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44930;
    wire N__44929;
    wire N__44926;
    wire N__44921;
    wire N__44916;
    wire N__44915;
    wire N__44914;
    wire N__44911;
    wire N__44908;
    wire N__44903;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44886;
    wire N__44885;
    wire N__44884;
    wire N__44881;
    wire N__44878;
    wire N__44875;
    wire N__44872;
    wire N__44871;
    wire N__44868;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44852;
    wire N__44847;
    wire N__44844;
    wire N__44843;
    wire N__44842;
    wire N__44839;
    wire N__44834;
    wire N__44831;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44821;
    wire N__44818;
    wire N__44815;
    wire N__44808;
    wire N__44807;
    wire N__44806;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44796;
    wire N__44793;
    wire N__44790;
    wire N__44787;
    wire N__44784;
    wire N__44779;
    wire N__44774;
    wire N__44769;
    wire N__44768;
    wire N__44767;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44755;
    wire N__44754;
    wire N__44751;
    wire N__44746;
    wire N__44743;
    wire N__44740;
    wire N__44735;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44721;
    wire N__44718;
    wire N__44717;
    wire N__44716;
    wire N__44713;
    wire N__44710;
    wire N__44707;
    wire N__44706;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44692;
    wire N__44689;
    wire N__44686;
    wire N__44683;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44643;
    wire N__44642;
    wire N__44639;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44622;
    wire N__44621;
    wire N__44618;
    wire N__44617;
    wire N__44616;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44601;
    wire N__44598;
    wire N__44591;
    wire N__44586;
    wire N__44583;
    wire N__44580;
    wire N__44577;
    wire N__44574;
    wire N__44571;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44563;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44547;
    wire N__44544;
    wire N__44543;
    wire N__44540;
    wire N__44537;
    wire N__44536;
    wire N__44531;
    wire N__44528;
    wire N__44525;
    wire N__44520;
    wire N__44517;
    wire N__44516;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44502;
    wire N__44499;
    wire N__44498;
    wire N__44497;
    wire N__44496;
    wire N__44495;
    wire N__44494;
    wire N__44493;
    wire N__44492;
    wire N__44491;
    wire N__44490;
    wire N__44489;
    wire N__44488;
    wire N__44487;
    wire N__44486;
    wire N__44485;
    wire N__44484;
    wire N__44483;
    wire N__44482;
    wire N__44481;
    wire N__44480;
    wire N__44479;
    wire N__44478;
    wire N__44477;
    wire N__44476;
    wire N__44475;
    wire N__44474;
    wire N__44473;
    wire N__44472;
    wire N__44471;
    wire N__44470;
    wire N__44463;
    wire N__44454;
    wire N__44445;
    wire N__44436;
    wire N__44427;
    wire N__44420;
    wire N__44411;
    wire N__44402;
    wire N__44393;
    wire N__44382;
    wire N__44379;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44364;
    wire N__44363;
    wire N__44360;
    wire N__44357;
    wire N__44356;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44343;
    wire N__44338;
    wire N__44333;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44321;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44308;
    wire N__44305;
    wire N__44298;
    wire N__44297;
    wire N__44296;
    wire N__44293;
    wire N__44290;
    wire N__44287;
    wire N__44286;
    wire N__44283;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44269;
    wire N__44266;
    wire N__44259;
    wire N__44256;
    wire N__44255;
    wire N__44252;
    wire N__44251;
    wire N__44248;
    wire N__44245;
    wire N__44242;
    wire N__44235;
    wire N__44234;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44218;
    wire N__44213;
    wire N__44210;
    wire N__44205;
    wire N__44202;
    wire N__44201;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44185;
    wire N__44178;
    wire N__44175;
    wire N__44174;
    wire N__44171;
    wire N__44168;
    wire N__44167;
    wire N__44162;
    wire N__44159;
    wire N__44156;
    wire N__44151;
    wire N__44148;
    wire N__44147;
    wire N__44144;
    wire N__44141;
    wire N__44140;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44124;
    wire N__44121;
    wire N__44120;
    wire N__44119;
    wire N__44114;
    wire N__44111;
    wire N__44108;
    wire N__44103;
    wire N__44100;
    wire N__44097;
    wire N__44096;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44081;
    wire N__44076;
    wire N__44073;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44065;
    wire N__44060;
    wire N__44057;
    wire N__44054;
    wire N__44049;
    wire N__44046;
    wire N__44045;
    wire N__44044;
    wire N__44039;
    wire N__44036;
    wire N__44033;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44014;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__43998;
    wire N__43995;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43975;
    wire N__43972;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43955;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43945;
    wire N__43942;
    wire N__43939;
    wire N__43932;
    wire N__43929;
    wire N__43928;
    wire N__43927;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43911;
    wire N__43908;
    wire N__43907;
    wire N__43902;
    wire N__43901;
    wire N__43898;
    wire N__43895;
    wire N__43892;
    wire N__43887;
    wire N__43884;
    wire N__43883;
    wire N__43880;
    wire N__43879;
    wire N__43876;
    wire N__43873;
    wire N__43870;
    wire N__43865;
    wire N__43860;
    wire N__43857;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43845;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43835;
    wire N__43830;
    wire N__43827;
    wire N__43826;
    wire N__43823;
    wire N__43820;
    wire N__43815;
    wire N__43814;
    wire N__43811;
    wire N__43808;
    wire N__43805;
    wire N__43800;
    wire N__43797;
    wire N__43796;
    wire N__43791;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43781;
    wire N__43776;
    wire N__43773;
    wire N__43770;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43762;
    wire N__43757;
    wire N__43754;
    wire N__43751;
    wire N__43746;
    wire N__43743;
    wire N__43742;
    wire N__43739;
    wire N__43736;
    wire N__43733;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43718;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43706;
    wire N__43703;
    wire N__43702;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43683;
    wire N__43680;
    wire N__43679;
    wire N__43676;
    wire N__43673;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43658;
    wire N__43653;
    wire N__43650;
    wire N__43649;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43639;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43623;
    wire N__43620;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43608;
    wire N__43607;
    wire N__43604;
    wire N__43601;
    wire N__43598;
    wire N__43593;
    wire N__43590;
    wire N__43589;
    wire N__43586;
    wire N__43583;
    wire N__43578;
    wire N__43577;
    wire N__43574;
    wire N__43571;
    wire N__43568;
    wire N__43563;
    wire N__43560;
    wire N__43559;
    wire N__43554;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43525;
    wire N__43520;
    wire N__43517;
    wire N__43514;
    wire N__43509;
    wire N__43506;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43492;
    wire N__43487;
    wire N__43484;
    wire N__43481;
    wire N__43476;
    wire N__43473;
    wire N__43472;
    wire N__43471;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43452;
    wire N__43449;
    wire N__43446;
    wire N__43443;
    wire N__43440;
    wire N__43431;
    wire N__43428;
    wire N__43427;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43416;
    wire N__43413;
    wire N__43408;
    wire N__43405;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43391;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43376;
    wire N__43373;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43363;
    wire N__43356;
    wire N__43353;
    wire N__43352;
    wire N__43347;
    wire N__43346;
    wire N__43343;
    wire N__43340;
    wire N__43335;
    wire N__43334;
    wire N__43331;
    wire N__43328;
    wire N__43323;
    wire N__43320;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43312;
    wire N__43307;
    wire N__43304;
    wire N__43303;
    wire N__43298;
    wire N__43295;
    wire N__43292;
    wire N__43289;
    wire N__43284;
    wire N__43281;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43264;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43254;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43236;
    wire N__43233;
    wire N__43232;
    wire N__43231;
    wire N__43230;
    wire N__43229;
    wire N__43228;
    wire N__43227;
    wire N__43226;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43197;
    wire N__43194;
    wire N__43193;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43166;
    wire N__43163;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43143;
    wire N__43140;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43132;
    wire N__43129;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43115;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43089;
    wire N__43088;
    wire N__43087;
    wire N__43084;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43070;
    wire N__43069;
    wire N__43066;
    wire N__43063;
    wire N__43060;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43046;
    wire N__43043;
    wire N__43042;
    wire N__43039;
    wire N__43036;
    wire N__43033;
    wire N__43030;
    wire N__43029;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43011;
    wire N__43008;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42981;
    wire N__42980;
    wire N__42977;
    wire N__42974;
    wire N__42969;
    wire N__42966;
    wire N__42965;
    wire N__42960;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42948;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42936;
    wire N__42933;
    wire N__42932;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42922;
    wire N__42917;
    wire N__42914;
    wire N__42913;
    wire N__42910;
    wire N__42907;
    wire N__42904;
    wire N__42897;
    wire N__42894;
    wire N__42893;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42880;
    wire N__42875;
    wire N__42874;
    wire N__42869;
    wire N__42866;
    wire N__42861;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42851;
    wire N__42848;
    wire N__42845;
    wire N__42842;
    wire N__42839;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42826;
    wire N__42821;
    wire N__42820;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42804;
    wire N__42801;
    wire N__42800;
    wire N__42797;
    wire N__42796;
    wire N__42793;
    wire N__42790;
    wire N__42787;
    wire N__42784;
    wire N__42781;
    wire N__42778;
    wire N__42777;
    wire N__42774;
    wire N__42769;
    wire N__42766;
    wire N__42759;
    wire N__42756;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42743;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42732;
    wire N__42725;
    wire N__42722;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42710;
    wire N__42709;
    wire N__42706;
    wire N__42701;
    wire N__42698;
    wire N__42695;
    wire N__42694;
    wire N__42691;
    wire N__42688;
    wire N__42685;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42671;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42658;
    wire N__42655;
    wire N__42652;
    wire N__42651;
    wire N__42648;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42631;
    wire N__42624;
    wire N__42621;
    wire N__42620;
    wire N__42617;
    wire N__42614;
    wire N__42613;
    wire N__42608;
    wire N__42605;
    wire N__42604;
    wire N__42599;
    wire N__42596;
    wire N__42593;
    wire N__42590;
    wire N__42585;
    wire N__42582;
    wire N__42581;
    wire N__42578;
    wire N__42577;
    wire N__42576;
    wire N__42573;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42557;
    wire N__42554;
    wire N__42551;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42489;
    wire N__42488;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42473;
    wire N__42472;
    wire N__42469;
    wire N__42466;
    wire N__42463;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42449;
    wire N__42446;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42431;
    wire N__42428;
    wire N__42427;
    wire N__42424;
    wire N__42421;
    wire N__42418;
    wire N__42411;
    wire N__42408;
    wire N__42407;
    wire N__42404;
    wire N__42401;
    wire N__42400;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42382;
    wire N__42379;
    wire N__42374;
    wire N__42371;
    wire N__42368;
    wire N__42363;
    wire N__42360;
    wire N__42359;
    wire N__42356;
    wire N__42353;
    wire N__42350;
    wire N__42347;
    wire N__42346;
    wire N__42345;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42296;
    wire N__42293;
    wire N__42290;
    wire N__42285;
    wire N__42284;
    wire N__42283;
    wire N__42278;
    wire N__42277;
    wire N__42274;
    wire N__42271;
    wire N__42268;
    wire N__42263;
    wire N__42260;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42242;
    wire N__42239;
    wire N__42236;
    wire N__42231;
    wire N__42230;
    wire N__42229;
    wire N__42226;
    wire N__42223;
    wire N__42220;
    wire N__42213;
    wire N__42212;
    wire N__42209;
    wire N__42206;
    wire N__42203;
    wire N__42200;
    wire N__42195;
    wire N__42192;
    wire N__42191;
    wire N__42190;
    wire N__42187;
    wire N__42184;
    wire N__42181;
    wire N__42174;
    wire N__42171;
    wire N__42168;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42150;
    wire N__42147;
    wire N__42144;
    wire N__42141;
    wire N__42138;
    wire N__42135;
    wire N__42132;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42122;
    wire N__42121;
    wire N__42120;
    wire N__42119;
    wire N__42118;
    wire N__42117;
    wire N__42116;
    wire N__42115;
    wire N__42114;
    wire N__42113;
    wire N__42112;
    wire N__42111;
    wire N__42110;
    wire N__42109;
    wire N__42108;
    wire N__42107;
    wire N__42106;
    wire N__42105;
    wire N__42104;
    wire N__42103;
    wire N__42102;
    wire N__42101;
    wire N__42100;
    wire N__42099;
    wire N__42098;
    wire N__42097;
    wire N__42096;
    wire N__42095;
    wire N__42094;
    wire N__42093;
    wire N__42092;
    wire N__42089;
    wire N__42086;
    wire N__42079;
    wire N__42070;
    wire N__42061;
    wire N__42052;
    wire N__42043;
    wire N__42034;
    wire N__42027;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42007;
    wire N__42002;
    wire N__41997;
    wire N__41992;
    wire N__41989;
    wire N__41984;
    wire N__41981;
    wire N__41978;
    wire N__41975;
    wire N__41970;
    wire N__41967;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41951;
    wire N__41948;
    wire N__41945;
    wire N__41944;
    wire N__41941;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41927;
    wire N__41924;
    wire N__41921;
    wire N__41918;
    wire N__41915;
    wire N__41912;
    wire N__41909;
    wire N__41904;
    wire N__41901;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41883;
    wire N__41882;
    wire N__41879;
    wire N__41876;
    wire N__41871;
    wire N__41868;
    wire N__41867;
    wire N__41864;
    wire N__41861;
    wire N__41858;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41841;
    wire N__41838;
    wire N__41835;
    wire N__41834;
    wire N__41833;
    wire N__41832;
    wire N__41829;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41812;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41798;
    wire N__41795;
    wire N__41792;
    wire N__41787;
    wire N__41786;
    wire N__41785;
    wire N__41778;
    wire N__41775;
    wire N__41774;
    wire N__41773;
    wire N__41772;
    wire N__41769;
    wire N__41762;
    wire N__41757;
    wire N__41756;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41748;
    wire N__41745;
    wire N__41738;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41723;
    wire N__41720;
    wire N__41719;
    wire N__41712;
    wire N__41709;
    wire N__41708;
    wire N__41707;
    wire N__41704;
    wire N__41699;
    wire N__41698;
    wire N__41693;
    wire N__41690;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41678;
    wire N__41675;
    wire N__41672;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41657;
    wire N__41656;
    wire N__41651;
    wire N__41648;
    wire N__41645;
    wire N__41640;
    wire N__41637;
    wire N__41634;
    wire N__41633;
    wire N__41632;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41616;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41577;
    wire N__41574;
    wire N__41573;
    wire N__41570;
    wire N__41567;
    wire N__41562;
    wire N__41559;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41547;
    wire N__41544;
    wire N__41543;
    wire N__41542;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41526;
    wire N__41523;
    wire N__41522;
    wire N__41519;
    wire N__41514;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41504;
    wire N__41499;
    wire N__41496;
    wire N__41495;
    wire N__41494;
    wire N__41489;
    wire N__41486;
    wire N__41483;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41471;
    wire N__41470;
    wire N__41465;
    wire N__41462;
    wire N__41459;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41433;
    wire N__41430;
    wire N__41427;
    wire N__41426;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41412;
    wire N__41409;
    wire N__41408;
    wire N__41405;
    wire N__41402;
    wire N__41397;
    wire N__41394;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41382;
    wire N__41379;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41364;
    wire N__41361;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41349;
    wire N__41346;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41334;
    wire N__41331;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41310;
    wire N__41307;
    wire N__41306;
    wire N__41303;
    wire N__41302;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41290;
    wire N__41283;
    wire N__41282;
    wire N__41281;
    wire N__41280;
    wire N__41279;
    wire N__41274;
    wire N__41271;
    wire N__41266;
    wire N__41259;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41247;
    wire N__41244;
    wire N__41243;
    wire N__41242;
    wire N__41239;
    wire N__41236;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41212;
    wire N__41209;
    wire N__41206;
    wire N__41203;
    wire N__41196;
    wire N__41193;
    wire N__41192;
    wire N__41191;
    wire N__41190;
    wire N__41189;
    wire N__41188;
    wire N__41187;
    wire N__41186;
    wire N__41185;
    wire N__41184;
    wire N__41183;
    wire N__41182;
    wire N__41181;
    wire N__41180;
    wire N__41179;
    wire N__41178;
    wire N__41177;
    wire N__41176;
    wire N__41175;
    wire N__41174;
    wire N__41173;
    wire N__41172;
    wire N__41171;
    wire N__41170;
    wire N__41169;
    wire N__41168;
    wire N__41167;
    wire N__41166;
    wire N__41165;
    wire N__41164;
    wire N__41163;
    wire N__41162;
    wire N__41161;
    wire N__41160;
    wire N__41159;
    wire N__41156;
    wire N__41147;
    wire N__41144;
    wire N__41143;
    wire N__41142;
    wire N__41139;
    wire N__41138;
    wire N__41137;
    wire N__41136;
    wire N__41135;
    wire N__41134;
    wire N__41133;
    wire N__41132;
    wire N__41129;
    wire N__41128;
    wire N__41127;
    wire N__41126;
    wire N__41125;
    wire N__41124;
    wire N__41123;
    wire N__41122;
    wire N__41121;
    wire N__41120;
    wire N__41119;
    wire N__41116;
    wire N__41115;
    wire N__41112;
    wire N__41111;
    wire N__41110;
    wire N__41109;
    wire N__41106;
    wire N__41105;
    wire N__41104;
    wire N__41099;
    wire N__41098;
    wire N__41097;
    wire N__41096;
    wire N__41095;
    wire N__41094;
    wire N__41093;
    wire N__41092;
    wire N__41087;
    wire N__41078;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41060;
    wire N__41057;
    wire N__41050;
    wire N__41045;
    wire N__41038;
    wire N__41031;
    wire N__41024;
    wire N__41021;
    wire N__41018;
    wire N__41011;
    wire N__41006;
    wire N__41003;
    wire N__41002;
    wire N__41001;
    wire N__41000;
    wire N__40999;
    wire N__40998;
    wire N__40997;
    wire N__40996;
    wire N__40995;
    wire N__40994;
    wire N__40993;
    wire N__40992;
    wire N__40991;
    wire N__40990;
    wire N__40973;
    wire N__40964;
    wire N__40961;
    wire N__40958;
    wire N__40957;
    wire N__40956;
    wire N__40955;
    wire N__40954;
    wire N__40953;
    wire N__40952;
    wire N__40951;
    wire N__40950;
    wire N__40949;
    wire N__40948;
    wire N__40947;
    wire N__40946;
    wire N__40941;
    wire N__40938;
    wire N__40933;
    wire N__40930;
    wire N__40919;
    wire N__40914;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40886;
    wire N__40881;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40857;
    wire N__40844;
    wire N__40837;
    wire N__40828;
    wire N__40821;
    wire N__40814;
    wire N__40807;
    wire N__40798;
    wire N__40789;
    wire N__40778;
    wire N__40755;
    wire N__40752;
    wire N__40751;
    wire N__40748;
    wire N__40745;
    wire N__40742;
    wire N__40739;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40716;
    wire N__40715;
    wire N__40712;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40682;
    wire N__40679;
    wire N__40676;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40662;
    wire N__40659;
    wire N__40658;
    wire N__40655;
    wire N__40652;
    wire N__40647;
    wire N__40644;
    wire N__40643;
    wire N__40640;
    wire N__40637;
    wire N__40632;
    wire N__40629;
    wire N__40628;
    wire N__40627;
    wire N__40626;
    wire N__40625;
    wire N__40622;
    wire N__40621;
    wire N__40618;
    wire N__40617;
    wire N__40616;
    wire N__40615;
    wire N__40614;
    wire N__40613;
    wire N__40612;
    wire N__40611;
    wire N__40610;
    wire N__40609;
    wire N__40608;
    wire N__40607;
    wire N__40606;
    wire N__40605;
    wire N__40604;
    wire N__40603;
    wire N__40602;
    wire N__40601;
    wire N__40600;
    wire N__40599;
    wire N__40598;
    wire N__40597;
    wire N__40596;
    wire N__40595;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40587;
    wire N__40586;
    wire N__40585;
    wire N__40584;
    wire N__40583;
    wire N__40582;
    wire N__40581;
    wire N__40580;
    wire N__40579;
    wire N__40578;
    wire N__40577;
    wire N__40576;
    wire N__40575;
    wire N__40574;
    wire N__40573;
    wire N__40572;
    wire N__40571;
    wire N__40570;
    wire N__40567;
    wire N__40566;
    wire N__40565;
    wire N__40564;
    wire N__40561;
    wire N__40544;
    wire N__40531;
    wire N__40528;
    wire N__40519;
    wire N__40512;
    wire N__40507;
    wire N__40502;
    wire N__40487;
    wire N__40486;
    wire N__40485;
    wire N__40484;
    wire N__40483;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40466;
    wire N__40453;
    wire N__40452;
    wire N__40451;
    wire N__40450;
    wire N__40449;
    wire N__40448;
    wire N__40447;
    wire N__40446;
    wire N__40445;
    wire N__40444;
    wire N__40443;
    wire N__40442;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40428;
    wire N__40423;
    wire N__40420;
    wire N__40417;
    wire N__40412;
    wire N__40407;
    wire N__40404;
    wire N__40393;
    wire N__40388;
    wire N__40381;
    wire N__40364;
    wire N__40363;
    wire N__40362;
    wire N__40361;
    wire N__40358;
    wire N__40351;
    wire N__40344;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40326;
    wire N__40319;
    wire N__40312;
    wire N__40293;
    wire N__40292;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40279;
    wire N__40272;
    wire N__40271;
    wire N__40270;
    wire N__40269;
    wire N__40268;
    wire N__40267;
    wire N__40266;
    wire N__40265;
    wire N__40264;
    wire N__40263;
    wire N__40262;
    wire N__40261;
    wire N__40260;
    wire N__40257;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40247;
    wire N__40246;
    wire N__40245;
    wire N__40242;
    wire N__40239;
    wire N__40238;
    wire N__40237;
    wire N__40236;
    wire N__40235;
    wire N__40234;
    wire N__40233;
    wire N__40232;
    wire N__40231;
    wire N__40230;
    wire N__40229;
    wire N__40228;
    wire N__40225;
    wire N__40218;
    wire N__40209;
    wire N__40208;
    wire N__40205;
    wire N__40204;
    wire N__40203;
    wire N__40202;
    wire N__40201;
    wire N__40200;
    wire N__40199;
    wire N__40198;
    wire N__40197;
    wire N__40196;
    wire N__40195;
    wire N__40192;
    wire N__40187;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40175;
    wire N__40174;
    wire N__40171;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40151;
    wire N__40150;
    wire N__40147;
    wire N__40146;
    wire N__40145;
    wire N__40144;
    wire N__40143;
    wire N__40142;
    wire N__40141;
    wire N__40140;
    wire N__40139;
    wire N__40138;
    wire N__40137;
    wire N__40136;
    wire N__40135;
    wire N__40134;
    wire N__40133;
    wire N__40130;
    wire N__40129;
    wire N__40128;
    wire N__40127;
    wire N__40126;
    wire N__40125;
    wire N__40122;
    wire N__40121;
    wire N__40120;
    wire N__40115;
    wire N__40114;
    wire N__40113;
    wire N__40112;
    wire N__40111;
    wire N__40106;
    wire N__40101;
    wire N__40086;
    wire N__40079;
    wire N__40076;
    wire N__40073;
    wire N__40066;
    wire N__40061;
    wire N__40052;
    wire N__40043;
    wire N__40040;
    wire N__40035;
    wire N__40034;
    wire N__40033;
    wire N__40030;
    wire N__40029;
    wire N__40026;
    wire N__40025;
    wire N__40022;
    wire N__40021;
    wire N__40020;
    wire N__40017;
    wire N__40016;
    wire N__40013;
    wire N__40012;
    wire N__40009;
    wire N__40008;
    wire N__40007;
    wire N__40004;
    wire N__40003;
    wire N__40000;
    wire N__39999;
    wire N__39996;
    wire N__39995;
    wire N__39992;
    wire N__39989;
    wire N__39988;
    wire N__39985;
    wire N__39984;
    wire N__39981;
    wire N__39980;
    wire N__39977;
    wire N__39976;
    wire N__39975;
    wire N__39974;
    wire N__39973;
    wire N__39972;
    wire N__39971;
    wire N__39970;
    wire N__39969;
    wire N__39968;
    wire N__39967;
    wire N__39966;
    wire N__39965;
    wire N__39962;
    wire N__39959;
    wire N__39958;
    wire N__39957;
    wire N__39956;
    wire N__39955;
    wire N__39954;
    wire N__39939;
    wire N__39936;
    wire N__39927;
    wire N__39918;
    wire N__39901;
    wire N__39884;
    wire N__39869;
    wire N__39852;
    wire N__39835;
    wire N__39832;
    wire N__39831;
    wire N__39828;
    wire N__39827;
    wire N__39824;
    wire N__39823;
    wire N__39820;
    wire N__39819;
    wire N__39816;
    wire N__39815;
    wire N__39812;
    wire N__39811;
    wire N__39808;
    wire N__39807;
    wire N__39804;
    wire N__39803;
    wire N__39802;
    wire N__39801;
    wire N__39800;
    wire N__39799;
    wire N__39796;
    wire N__39795;
    wire N__39792;
    wire N__39791;
    wire N__39788;
    wire N__39787;
    wire N__39786;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39768;
    wire N__39765;
    wire N__39758;
    wire N__39747;
    wire N__39730;
    wire N__39713;
    wire N__39706;
    wire N__39693;
    wire N__39686;
    wire N__39663;
    wire N__39660;
    wire N__39657;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39636;
    wire N__39633;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39603;
    wire N__39600;
    wire N__39599;
    wire N__39596;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39576;
    wire N__39575;
    wire N__39572;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39537;
    wire N__39534;
    wire N__39531;
    wire N__39528;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39490;
    wire N__39487;
    wire N__39484;
    wire N__39481;
    wire N__39480;
    wire N__39477;
    wire N__39472;
    wire N__39469;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39453;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39445;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39437;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39411;
    wire N__39408;
    wire N__39407;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39365;
    wire N__39364;
    wire N__39361;
    wire N__39358;
    wire N__39355;
    wire N__39350;
    wire N__39345;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39272;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39258;
    wire N__39257;
    wire N__39254;
    wire N__39251;
    wire N__39248;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39233;
    wire N__39232;
    wire N__39225;
    wire N__39224;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39210;
    wire N__39207;
    wire N__39206;
    wire N__39203;
    wire N__39200;
    wire N__39197;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39185;
    wire N__39184;
    wire N__39179;
    wire N__39176;
    wire N__39173;
    wire N__39168;
    wire N__39165;
    wire N__39164;
    wire N__39163;
    wire N__39158;
    wire N__39155;
    wire N__39152;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39137;
    wire N__39134;
    wire N__39133;
    wire N__39128;
    wire N__39125;
    wire N__39122;
    wire N__39117;
    wire N__39114;
    wire N__39113;
    wire N__39112;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39089;
    wire N__39084;
    wire N__39083;
    wire N__39080;
    wire N__39077;
    wire N__39074;
    wire N__39069;
    wire N__39066;
    wire N__39065;
    wire N__39060;
    wire N__39059;
    wire N__39056;
    wire N__39053;
    wire N__39050;
    wire N__39045;
    wire N__39042;
    wire N__39041;
    wire N__39038;
    wire N__39035;
    wire N__39032;
    wire N__39027;
    wire N__39024;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39009;
    wire N__39006;
    wire N__39005;
    wire N__39002;
    wire N__38999;
    wire N__38996;
    wire N__38991;
    wire N__38988;
    wire N__38987;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38973;
    wire N__38970;
    wire N__38969;
    wire N__38966;
    wire N__38963;
    wire N__38960;
    wire N__38955;
    wire N__38952;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38937;
    wire N__38934;
    wire N__38933;
    wire N__38930;
    wire N__38927;
    wire N__38924;
    wire N__38919;
    wire N__38916;
    wire N__38915;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38892;
    wire N__38889;
    wire N__38886;
    wire N__38883;
    wire N__38882;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38855;
    wire N__38854;
    wire N__38851;
    wire N__38848;
    wire N__38845;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38830;
    wire N__38823;
    wire N__38822;
    wire N__38819;
    wire N__38816;
    wire N__38813;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38775;
    wire N__38772;
    wire N__38771;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38757;
    wire N__38754;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38456;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38448;
    wire N__38443;
    wire N__38438;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38417;
    wire N__38414;
    wire N__38411;
    wire N__38406;
    wire N__38403;
    wire N__38402;
    wire N__38399;
    wire N__38396;
    wire N__38391;
    wire N__38390;
    wire N__38387;
    wire N__38386;
    wire N__38385;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38367;
    wire N__38366;
    wire N__38363;
    wire N__38362;
    wire N__38361;
    wire N__38360;
    wire N__38355;
    wire N__38352;
    wire N__38347;
    wire N__38340;
    wire N__38337;
    wire N__38336;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38324;
    wire N__38319;
    wire N__38316;
    wire N__38315;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38276;
    wire N__38271;
    wire N__38270;
    wire N__38267;
    wire N__38264;
    wire N__38261;
    wire N__38256;
    wire N__38255;
    wire N__38252;
    wire N__38249;
    wire N__38248;
    wire N__38247;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38226;
    wire N__38225;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38213;
    wire N__38212;
    wire N__38207;
    wire N__38204;
    wire N__38199;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38187;
    wire N__38184;
    wire N__38181;
    wire N__38180;
    wire N__38177;
    wire N__38174;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38133;
    wire N__38132;
    wire N__38131;
    wire N__38128;
    wire N__38123;
    wire N__38122;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38106;
    wire N__38105;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38072;
    wire N__38069;
    wire N__38064;
    wire N__38063;
    wire N__38060;
    wire N__38057;
    wire N__38054;
    wire N__38051;
    wire N__38046;
    wire N__38043;
    wire N__38040;
    wire N__38039;
    wire N__38038;
    wire N__38037;
    wire N__38036;
    wire N__38035;
    wire N__38034;
    wire N__38019;
    wire N__38018;
    wire N__38017;
    wire N__38016;
    wire N__38015;
    wire N__38014;
    wire N__38013;
    wire N__38012;
    wire N__38011;
    wire N__38010;
    wire N__38009;
    wire N__38008;
    wire N__38007;
    wire N__38006;
    wire N__38005;
    wire N__38004;
    wire N__38003;
    wire N__38002;
    wire N__37999;
    wire N__37994;
    wire N__37991;
    wire N__37980;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37958;
    wire N__37957;
    wire N__37952;
    wire N__37947;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37917;
    wire N__37916;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37901;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37874;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37859;
    wire N__37854;
    wire N__37851;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37829;
    wire N__37828;
    wire N__37825;
    wire N__37822;
    wire N__37819;
    wire N__37814;
    wire N__37809;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37776;
    wire N__37775;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37765;
    wire N__37762;
    wire N__37759;
    wire N__37752;
    wire N__37749;
    wire N__37746;
    wire N__37743;
    wire N__37742;
    wire N__37741;
    wire N__37738;
    wire N__37735;
    wire N__37730;
    wire N__37727;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37712;
    wire N__37709;
    wire N__37708;
    wire N__37705;
    wire N__37702;
    wire N__37699;
    wire N__37696;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37682;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37662;
    wire N__37659;
    wire N__37656;
    wire N__37655;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37616;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37581;
    wire N__37578;
    wire N__37575;
    wire N__37574;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37559;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37537;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37499;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37487;
    wire N__37484;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37472;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37462;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37423;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37383;
    wire N__37380;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37302;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37248;
    wire N__37245;
    wire N__37242;
    wire N__37239;
    wire N__37236;
    wire N__37235;
    wire N__37234;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37183;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37167;
    wire N__37164;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37152;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37119;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37093;
    wire N__37090;
    wire N__37085;
    wire N__37080;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37054;
    wire N__37049;
    wire N__37046;
    wire N__37041;
    wire N__37038;
    wire N__37035;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36924;
    wire N__36921;
    wire N__36920;
    wire N__36917;
    wire N__36916;
    wire N__36913;
    wire N__36912;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36892;
    wire N__36885;
    wire N__36882;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36852;
    wire N__36849;
    wire N__36848;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36819;
    wire N__36816;
    wire N__36815;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36786;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36774;
    wire N__36771;
    wire N__36768;
    wire N__36765;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36741;
    wire N__36738;
    wire N__36737;
    wire N__36736;
    wire N__36735;
    wire N__36730;
    wire N__36727;
    wire N__36724;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36698;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36666;
    wire N__36663;
    wire N__36662;
    wire N__36661;
    wire N__36658;
    wire N__36653;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36643;
    wire N__36640;
    wire N__36637;
    wire N__36634;
    wire N__36627;
    wire N__36626;
    wire N__36621;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36604;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36569;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36557;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36540;
    wire N__36539;
    wire N__36536;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36519;
    wire N__36516;
    wire N__36515;
    wire N__36514;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36502;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36488;
    wire N__36485;
    wire N__36484;
    wire N__36481;
    wire N__36478;
    wire N__36475;
    wire N__36468;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36460;
    wire N__36459;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36428;
    wire N__36425;
    wire N__36424;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36408;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36400;
    wire N__36399;
    wire N__36394;
    wire N__36389;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36371;
    wire N__36370;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36339;
    wire N__36336;
    wire N__36333;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36321;
    wire N__36320;
    wire N__36315;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36294;
    wire N__36293;
    wire N__36292;
    wire N__36289;
    wire N__36284;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36267;
    wire N__36264;
    wire N__36263;
    wire N__36258;
    wire N__36255;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36243;
    wire N__36240;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36211;
    wire N__36204;
    wire N__36203;
    wire N__36200;
    wire N__36197;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36154;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36120;
    wire N__36119;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36107;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36089;
    wire N__36088;
    wire N__36085;
    wire N__36082;
    wire N__36081;
    wire N__36080;
    wire N__36079;
    wire N__36078;
    wire N__36077;
    wire N__36076;
    wire N__36075;
    wire N__36070;
    wire N__36067;
    wire N__36052;
    wire N__36049;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36029;
    wire N__36026;
    wire N__36021;
    wire N__36020;
    wire N__36019;
    wire N__36018;
    wire N__36017;
    wire N__36016;
    wire N__36015;
    wire N__36014;
    wire N__36013;
    wire N__36012;
    wire N__36011;
    wire N__36010;
    wire N__36009;
    wire N__36008;
    wire N__36007;
    wire N__36006;
    wire N__36005;
    wire N__36004;
    wire N__36003;
    wire N__36002;
    wire N__36001;
    wire N__36000;
    wire N__35999;
    wire N__35998;
    wire N__35993;
    wire N__35986;
    wire N__35969;
    wire N__35954;
    wire N__35953;
    wire N__35952;
    wire N__35951;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35943;
    wire N__35940;
    wire N__35939;
    wire N__35936;
    wire N__35931;
    wire N__35926;
    wire N__35921;
    wire N__35906;
    wire N__35903;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35888;
    wire N__35885;
    wire N__35884;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35867;
    wire N__35862;
    wire N__35853;
    wire N__35852;
    wire N__35847;
    wire N__35846;
    wire N__35843;
    wire N__35842;
    wire N__35841;
    wire N__35840;
    wire N__35839;
    wire N__35838;
    wire N__35837;
    wire N__35836;
    wire N__35833;
    wire N__35830;
    wire N__35815;
    wire N__35812;
    wire N__35805;
    wire N__35802;
    wire N__35799;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35777;
    wire N__35774;
    wire N__35769;
    wire N__35766;
    wire N__35763;
    wire N__35760;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35739;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35731;
    wire N__35726;
    wire N__35723;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35709;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35691;
    wire N__35688;
    wire N__35685;
    wire N__35682;
    wire N__35679;
    wire N__35676;
    wire N__35675;
    wire N__35672;
    wire N__35671;
    wire N__35670;
    wire N__35669;
    wire N__35668;
    wire N__35665;
    wire N__35664;
    wire N__35663;
    wire N__35662;
    wire N__35661;
    wire N__35660;
    wire N__35659;
    wire N__35658;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35646;
    wire N__35643;
    wire N__35642;
    wire N__35641;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35627;
    wire N__35618;
    wire N__35611;
    wire N__35608;
    wire N__35607;
    wire N__35604;
    wire N__35601;
    wire N__35598;
    wire N__35597;
    wire N__35596;
    wire N__35595;
    wire N__35594;
    wire N__35593;
    wire N__35592;
    wire N__35591;
    wire N__35590;
    wire N__35589;
    wire N__35588;
    wire N__35587;
    wire N__35586;
    wire N__35585;
    wire N__35584;
    wire N__35583;
    wire N__35582;
    wire N__35581;
    wire N__35572;
    wire N__35569;
    wire N__35566;
    wire N__35563;
    wire N__35560;
    wire N__35555;
    wire N__35548;
    wire N__35539;
    wire N__35538;
    wire N__35537;
    wire N__35534;
    wire N__35533;
    wire N__35530;
    wire N__35529;
    wire N__35526;
    wire N__35525;
    wire N__35524;
    wire N__35521;
    wire N__35520;
    wire N__35517;
    wire N__35516;
    wire N__35513;
    wire N__35512;
    wire N__35509;
    wire N__35508;
    wire N__35507;
    wire N__35506;
    wire N__35505;
    wire N__35504;
    wire N__35503;
    wire N__35502;
    wire N__35501;
    wire N__35500;
    wire N__35495;
    wire N__35492;
    wire N__35489;
    wire N__35484;
    wire N__35481;
    wire N__35472;
    wire N__35471;
    wire N__35468;
    wire N__35467;
    wire N__35452;
    wire N__35435;
    wire N__35430;
    wire N__35427;
    wire N__35426;
    wire N__35423;
    wire N__35422;
    wire N__35419;
    wire N__35418;
    wire N__35415;
    wire N__35414;
    wire N__35413;
    wire N__35410;
    wire N__35409;
    wire N__35406;
    wire N__35405;
    wire N__35402;
    wire N__35401;
    wire N__35396;
    wire N__35393;
    wire N__35386;
    wire N__35379;
    wire N__35372;
    wire N__35355;
    wire N__35340;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35328;
    wire N__35321;
    wire N__35318;
    wire N__35313;
    wire N__35308;
    wire N__35301;
    wire N__35298;
    wire N__35297;
    wire N__35296;
    wire N__35291;
    wire N__35290;
    wire N__35289;
    wire N__35288;
    wire N__35287;
    wire N__35286;
    wire N__35285;
    wire N__35284;
    wire N__35283;
    wire N__35282;
    wire N__35279;
    wire N__35278;
    wire N__35277;
    wire N__35276;
    wire N__35273;
    wire N__35258;
    wire N__35253;
    wire N__35250;
    wire N__35243;
    wire N__35238;
    wire N__35235;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35219;
    wire N__35214;
    wire N__35211;
    wire N__35210;
    wire N__35209;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35197;
    wire N__35194;
    wire N__35187;
    wire N__35186;
    wire N__35183;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35166;
    wire N__35165;
    wire N__35162;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35145;
    wire N__35144;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35124;
    wire N__35123;
    wire N__35120;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35103;
    wire N__35102;
    wire N__35099;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35082;
    wire N__35081;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35061;
    wire N__35060;
    wire N__35059;
    wire N__35056;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35040;
    wire N__35037;
    wire N__35036;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35016;
    wire N__35013;
    wire N__35010;
    wire N__35009;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34989;
    wire N__34986;
    wire N__34985;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34965;
    wire N__34964;
    wire N__34963;
    wire N__34962;
    wire N__34961;
    wire N__34960;
    wire N__34959;
    wire N__34958;
    wire N__34957;
    wire N__34956;
    wire N__34947;
    wire N__34942;
    wire N__34933;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34757;
    wire N__34754;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34656;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34554;
    wire N__34551;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34349;
    wire N__34348;
    wire N__34347;
    wire N__34346;
    wire N__34345;
    wire N__34344;
    wire N__34343;
    wire N__34342;
    wire N__34341;
    wire N__34340;
    wire N__34339;
    wire N__34338;
    wire N__34337;
    wire N__34336;
    wire N__34335;
    wire N__34334;
    wire N__34333;
    wire N__34332;
    wire N__34331;
    wire N__34322;
    wire N__34313;
    wire N__34312;
    wire N__34311;
    wire N__34310;
    wire N__34309;
    wire N__34308;
    wire N__34307;
    wire N__34306;
    wire N__34305;
    wire N__34304;
    wire N__34303;
    wire N__34294;
    wire N__34285;
    wire N__34276;
    wire N__34271;
    wire N__34266;
    wire N__34257;
    wire N__34248;
    wire N__34245;
    wire N__34238;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34210;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34194;
    wire N__34191;
    wire N__34190;
    wire N__34189;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34173;
    wire N__34170;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34148;
    wire N__34143;
    wire N__34140;
    wire N__34139;
    wire N__34136;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34103;
    wire N__34100;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34083;
    wire N__34080;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34072;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34056;
    wire N__34053;
    wire N__34052;
    wire N__34051;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34035;
    wire N__34032;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33993;
    wire N__33992;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33939;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33931;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33915;
    wire N__33912;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33900;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33885;
    wire N__33882;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33860;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33846;
    wire N__33845;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33828;
    wire N__33825;
    wire N__33822;
    wire N__33819;
    wire N__33818;
    wire N__33815;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33798;
    wire N__33795;
    wire N__33794;
    wire N__33793;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33770;
    wire N__33769;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33753;
    wire N__33750;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33738;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33723;
    wire N__33720;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33712;
    wire N__33707;
    wire N__33704;
    wire N__33701;
    wire N__33696;
    wire N__33693;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33681;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33652;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33626;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33599;
    wire N__33596;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33579;
    wire N__33576;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33568;
    wire N__33563;
    wire N__33560;
    wire N__33557;
    wire N__33552;
    wire N__33549;
    wire N__33548;
    wire N__33547;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33531;
    wire N__33528;
    wire N__33527;
    wire N__33526;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33461;
    wire N__33458;
    wire N__33457;
    wire N__33454;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33433;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33407;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33380;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33365;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33353;
    wire N__33352;
    wire N__33347;
    wire N__33344;
    wire N__33341;
    wire N__33336;
    wire N__33333;
    wire N__33332;
    wire N__33331;
    wire N__33326;
    wire N__33323;
    wire N__33320;
    wire N__33315;
    wire N__33312;
    wire N__33309;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33155;
    wire N__33152;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33132;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33079;
    wire N__33078;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33041;
    wire N__33040;
    wire N__33039;
    wire N__33032;
    wire N__33029;
    wire N__33024;
    wire N__33021;
    wire N__33020;
    wire N__33019;
    wire N__33018;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32856;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32797;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32753;
    wire N__32750;
    wire N__32749;
    wire N__32746;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32731;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32715;
    wire N__32714;
    wire N__32713;
    wire N__32710;
    wire N__32705;
    wire N__32700;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32689;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32673;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32654;
    wire N__32653;
    wire N__32650;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32615;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32603;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32591;
    wire N__32590;
    wire N__32583;
    wire N__32580;
    wire N__32579;
    wire N__32578;
    wire N__32571;
    wire N__32568;
    wire N__32565;
    wire N__32562;
    wire N__32559;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32484;
    wire N__32481;
    wire N__32480;
    wire N__32479;
    wire N__32478;
    wire N__32477;
    wire N__32476;
    wire N__32475;
    wire N__32474;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32468;
    wire N__32467;
    wire N__32466;
    wire N__32465;
    wire N__32464;
    wire N__32463;
    wire N__32462;
    wire N__32461;
    wire N__32460;
    wire N__32459;
    wire N__32458;
    wire N__32457;
    wire N__32456;
    wire N__32455;
    wire N__32454;
    wire N__32453;
    wire N__32452;
    wire N__32451;
    wire N__32450;
    wire N__32449;
    wire N__32448;
    wire N__32447;
    wire N__32440;
    wire N__32431;
    wire N__32428;
    wire N__32425;
    wire N__32416;
    wire N__32407;
    wire N__32400;
    wire N__32391;
    wire N__32382;
    wire N__32373;
    wire N__32368;
    wire N__32365;
    wire N__32362;
    wire N__32357;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32319;
    wire N__32316;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32295;
    wire N__32294;
    wire N__32291;
    wire N__32290;
    wire N__32289;
    wire N__32280;
    wire N__32277;
    wire N__32276;
    wire N__32275;
    wire N__32274;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32250;
    wire N__32249;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32232;
    wire N__32229;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32217;
    wire N__32216;
    wire N__32215;
    wire N__32214;
    wire N__32211;
    wire N__32204;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32190;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32159;
    wire N__32158;
    wire N__32157;
    wire N__32154;
    wire N__32147;
    wire N__32142;
    wire N__32139;
    wire N__32138;
    wire N__32137;
    wire N__32134;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32112;
    wire N__32111;
    wire N__32108;
    wire N__32107;
    wire N__32106;
    wire N__32105;
    wire N__32102;
    wire N__32101;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32084;
    wire N__32083;
    wire N__32082;
    wire N__32081;
    wire N__32080;
    wire N__32079;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32071;
    wire N__32070;
    wire N__32069;
    wire N__32068;
    wire N__32067;
    wire N__32062;
    wire N__32057;
    wire N__32054;
    wire N__32053;
    wire N__32052;
    wire N__32051;
    wire N__32050;
    wire N__32049;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32029;
    wire N__32028;
    wire N__32027;
    wire N__32026;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32018;
    wire N__32017;
    wire N__32016;
    wire N__32015;
    wire N__32014;
    wire N__32011;
    wire N__32008;
    wire N__32001;
    wire N__31994;
    wire N__31985;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31968;
    wire N__31967;
    wire N__31966;
    wire N__31965;
    wire N__31964;
    wire N__31963;
    wire N__31962;
    wire N__31961;
    wire N__31960;
    wire N__31959;
    wire N__31958;
    wire N__31957;
    wire N__31956;
    wire N__31953;
    wire N__31944;
    wire N__31939;
    wire N__31936;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31913;
    wire N__31910;
    wire N__31907;
    wire N__31902;
    wire N__31899;
    wire N__31890;
    wire N__31881;
    wire N__31872;
    wire N__31865;
    wire N__31856;
    wire N__31851;
    wire N__31830;
    wire N__31827;
    wire N__31826;
    wire N__31823;
    wire N__31822;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31784;
    wire N__31783;
    wire N__31780;
    wire N__31775;
    wire N__31770;
    wire N__31769;
    wire N__31768;
    wire N__31761;
    wire N__31760;
    wire N__31759;
    wire N__31756;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31593;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31493;
    wire N__31492;
    wire N__31491;
    wire N__31484;
    wire N__31481;
    wire N__31478;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31466;
    wire N__31463;
    wire N__31462;
    wire N__31459;
    wire N__31452;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31437;
    wire N__31436;
    wire N__31433;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31370;
    wire N__31365;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31350;
    wire N__31347;
    wire N__31346;
    wire N__31341;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31319;
    wire N__31314;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31299;
    wire N__31296;
    wire N__31295;
    wire N__31294;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31278;
    wire N__31275;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31253;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31241;
    wire N__31238;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31208;
    wire N__31203;
    wire N__31202;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31188;
    wire N__31185;
    wire N__31184;
    wire N__31179;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31169;
    wire N__31164;
    wire N__31161;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31149;
    wire N__31146;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31134;
    wire N__31131;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31112;
    wire N__31107;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31092;
    wire N__31089;
    wire N__31088;
    wire N__31087;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31071;
    wire N__31068;
    wire N__31067;
    wire N__31062;
    wire N__31061;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31040;
    wire N__31035;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31020;
    wire N__31017;
    wire N__31016;
    wire N__31011;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30989;
    wire N__30984;
    wire N__30983;
    wire N__30980;
    wire N__30977;
    wire N__30974;
    wire N__30969;
    wire N__30966;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30954;
    wire N__30951;
    wire N__30950;
    wire N__30947;
    wire N__30944;
    wire N__30939;
    wire N__30936;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30924;
    wire N__30921;
    wire N__30920;
    wire N__30917;
    wire N__30914;
    wire N__30909;
    wire N__30906;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30894;
    wire N__30891;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30879;
    wire N__30876;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30864;
    wire N__30861;
    wire N__30860;
    wire N__30857;
    wire N__30854;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30758;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30740;
    wire N__30737;
    wire N__30736;
    wire N__30733;
    wire N__30730;
    wire N__30727;
    wire N__30720;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30684;
    wire N__30681;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30669;
    wire N__30666;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30620;
    wire N__30617;
    wire N__30614;
    wire N__30611;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30564;
    wire N__30561;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30419;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30356;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30342;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30282;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30221;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30152;
    wire N__30151;
    wire N__30150;
    wire N__30141;
    wire N__30138;
    wire N__30137;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30129;
    wire N__30128;
    wire N__30125;
    wire N__30116;
    wire N__30113;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30096;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29997;
    wire N__29994;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29936;
    wire N__29933;
    wire N__29932;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29895;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29885;
    wire N__29882;
    wire N__29881;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29869;
    wire N__29868;
    wire N__29867;
    wire N__29866;
    wire N__29863;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29843;
    wire N__29840;
    wire N__29835;
    wire N__29832;
    wire N__29831;
    wire N__29830;
    wire N__29829;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29780;
    wire N__29777;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29715;
    wire N__29714;
    wire N__29713;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29694;
    wire N__29693;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29681;
    wire N__29680;
    wire N__29677;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29637;
    wire N__29636;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29623;
    wire N__29620;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29588;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29097;
    wire N__29094;
    wire N__29091;
    wire N__29088;
    wire N__29085;
    wire N__29082;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29058;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28869;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28854;
    wire N__28851;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28799;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28773;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28676;
    wire N__28675;
    wire N__28674;
    wire N__28671;
    wire N__28664;
    wire N__28659;
    wire N__28658;
    wire N__28657;
    wire N__28650;
    wire N__28647;
    wire N__28646;
    wire N__28645;
    wire N__28642;
    wire N__28641;
    wire N__28638;
    wire N__28631;
    wire N__28626;
    wire N__28625;
    wire N__28622;
    wire N__28621;
    wire N__28618;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28604;
    wire N__28603;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28589;
    wire N__28586;
    wire N__28585;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28555;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28532;
    wire N__28531;
    wire N__28528;
    wire N__28523;
    wire N__28518;
    wire N__28515;
    wire N__28514;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28502;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28487;
    wire N__28486;
    wire N__28483;
    wire N__28478;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28445;
    wire N__28444;
    wire N__28441;
    wire N__28436;
    wire N__28431;
    wire N__28430;
    wire N__28429;
    wire N__28424;
    wire N__28421;
    wire N__28418;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28406;
    wire N__28405;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28389;
    wire N__28386;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28372;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28356;
    wire N__28353;
    wire N__28352;
    wire N__28349;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28326;
    wire N__28323;
    wire N__28322;
    wire N__28319;
    wire N__28318;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28295;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28280;
    wire N__28275;
    wire N__28272;
    wire N__28271;
    wire N__28270;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28254;
    wire N__28251;
    wire N__28250;
    wire N__28247;
    wire N__28246;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28230;
    wire N__28227;
    wire N__28226;
    wire N__28225;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28187;
    wire N__28186;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28170;
    wire N__28167;
    wire N__28166;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28154;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28142;
    wire N__28141;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27963;
    wire N__27960;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27914;
    wire N__27913;
    wire N__27912;
    wire N__27911;
    wire N__27910;
    wire N__27909;
    wire N__27908;
    wire N__27903;
    wire N__27896;
    wire N__27889;
    wire N__27886;
    wire N__27881;
    wire N__27878;
    wire N__27875;
    wire N__27870;
    wire N__27867;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27494;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27446;
    wire N__27443;
    wire N__27440;
    wire N__27435;
    wire N__27432;
    wire N__27431;
    wire N__27428;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27392;
    wire N__27389;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27372;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27333;
    wire N__27330;
    wire N__27329;
    wire N__27326;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27309;
    wire N__27308;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27230;
    wire N__27227;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27101;
    wire N__27098;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27081;
    wire N__27080;
    wire N__27079;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27038;
    wire N__27033;
    wire N__27030;
    wire N__27029;
    wire N__27024;
    wire N__27021;
    wire N__27020;
    wire N__27019;
    wire N__27018;
    wire N__27017;
    wire N__27016;
    wire N__27015;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26993;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26979;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26967;
    wire N__26966;
    wire N__26965;
    wire N__26964;
    wire N__26961;
    wire N__26954;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26912;
    wire N__26911;
    wire N__26910;
    wire N__26909;
    wire N__26908;
    wire N__26905;
    wire N__26904;
    wire N__26903;
    wire N__26902;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26886;
    wire N__26883;
    wire N__26878;
    wire N__26873;
    wire N__26870;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26854;
    wire N__26851;
    wire N__26844;
    wire N__26843;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26831;
    wire N__26828;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26811;
    wire N__26808;
    wire N__26807;
    wire N__26806;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26794;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26775;
    wire N__26772;
    wire N__26771;
    wire N__26766;
    wire N__26763;
    wire N__26762;
    wire N__26759;
    wire N__26758;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26725;
    wire N__26718;
    wire N__26717;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26694;
    wire N__26693;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26664;
    wire N__26663;
    wire N__26662;
    wire N__26661;
    wire N__26658;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26628;
    wire N__26625;
    wire N__26624;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26603;
    wire N__26600;
    wire N__26595;
    wire N__26594;
    wire N__26591;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26580;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26561;
    wire N__26556;
    wire N__26555;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26543;
    wire N__26540;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26523;
    wire N__26522;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26484;
    wire N__26475;
    wire N__26472;
    wire N__26471;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26459;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26443;
    wire N__26436;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26425;
    wire N__26424;
    wire N__26419;
    wire N__26414;
    wire N__26409;
    wire N__26406;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26394;
    wire N__26391;
    wire N__26390;
    wire N__26389;
    wire N__26388;
    wire N__26383;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26364;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26356;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26335;
    wire N__26332;
    wire N__26327;
    wire N__26324;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26312;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26289;
    wire N__26288;
    wire N__26287;
    wire N__26286;
    wire N__26283;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26261;
    wire N__26258;
    wire N__26253;
    wire N__26252;
    wire N__26247;
    wire N__26244;
    wire N__26243;
    wire N__26240;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26223;
    wire N__26222;
    wire N__26219;
    wire N__26218;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26195;
    wire N__26190;
    wire N__26187;
    wire N__26186;
    wire N__26181;
    wire N__26178;
    wire N__26177;
    wire N__26176;
    wire N__26171;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26142;
    wire N__26139;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26127;
    wire N__26124;
    wire N__26123;
    wire N__26118;
    wire N__26115;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26104;
    wire N__26103;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26085;
    wire N__26082;
    wire N__26081;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26058;
    wire N__26057;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26047;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26013;
    wire N__26012;
    wire N__26009;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25982;
    wire N__25981;
    wire N__25978;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25957;
    wire N__25954;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25907;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25886;
    wire N__25883;
    wire N__25878;
    wire N__25875;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25867;
    wire N__25866;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25850;
    wire N__25847;
    wire N__25842;
    wire N__25841;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25815;
    wire N__25812;
    wire N__25811;
    wire N__25806;
    wire N__25803;
    wire N__25802;
    wire N__25797;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25787;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25772;
    wire N__25767;
    wire N__25766;
    wire N__25763;
    wire N__25758;
    wire N__25755;
    wire N__25754;
    wire N__25749;
    wire N__25746;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25731;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25701;
    wire N__25700;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25670;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25658;
    wire N__25653;
    wire N__25650;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25547;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25472;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25459;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25436;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25424;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25398;
    wire N__25395;
    wire N__25394;
    wire N__25393;
    wire N__25390;
    wire N__25385;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25370;
    wire N__25367;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25349;
    wire N__25348;
    wire N__25347;
    wire N__25338;
    wire N__25337;
    wire N__25336;
    wire N__25335;
    wire N__25334;
    wire N__25333;
    wire N__25332;
    wire N__25331;
    wire N__25330;
    wire N__25329;
    wire N__25328;
    wire N__25327;
    wire N__25326;
    wire N__25325;
    wire N__25324;
    wire N__25323;
    wire N__25322;
    wire N__25321;
    wire N__25320;
    wire N__25319;
    wire N__25318;
    wire N__25317;
    wire N__25316;
    wire N__25315;
    wire N__25314;
    wire N__25313;
    wire N__25312;
    wire N__25309;
    wire N__25300;
    wire N__25295;
    wire N__25286;
    wire N__25277;
    wire N__25268;
    wire N__25259;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25234;
    wire N__25221;
    wire N__25220;
    wire N__25219;
    wire N__25218;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25176;
    wire N__25173;
    wire N__25164;
    wire N__25163;
    wire N__25160;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25143;
    wire N__25140;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25128;
    wire N__25127;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25110;
    wire N__25109;
    wire N__25104;
    wire N__25101;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25071;
    wire N__25070;
    wire N__25069;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25042;
    wire N__25039;
    wire N__25034;
    wire N__25029;
    wire N__25026;
    wire N__25025;
    wire N__25020;
    wire N__25017;
    wire N__25016;
    wire N__25015;
    wire N__25012;
    wire N__25011;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24992;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24969;
    wire N__24966;
    wire N__24965;
    wire N__24962;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24945;
    wire N__24944;
    wire N__24941;
    wire N__24940;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24916;
    wire N__24913;
    wire N__24906;
    wire N__24905;
    wire N__24902;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24885;
    wire N__24884;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24856;
    wire N__24851;
    wire N__24846;
    wire N__24843;
    wire N__24842;
    wire N__24841;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24819;
    wire N__24818;
    wire N__24815;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24805;
    wire N__24798;
    wire N__24797;
    wire N__24794;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24777;
    wire N__24776;
    wire N__24773;
    wire N__24772;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24733;
    wire N__24726;
    wire N__24723;
    wire N__24722;
    wire N__24719;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24709;
    wire N__24702;
    wire N__24701;
    wire N__24698;
    wire N__24697;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24669;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24661;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24649;
    wire N__24642;
    wire N__24639;
    wire N__24638;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24621;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24613;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24601;
    wire N__24598;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24582;
    wire N__24581;
    wire N__24578;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24561;
    wire N__24560;
    wire N__24557;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24547;
    wire N__24540;
    wire N__24537;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24508;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24494;
    wire N__24489;
    wire N__24486;
    wire N__24485;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24225;
    wire N__24222;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24195;
    wire N__24192;
    wire N__24189;
    wire N__24188;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24147;
    wire N__24144;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24092;
    wire N__24091;
    wire N__24088;
    wire N__24083;
    wire N__24078;
    wire N__24075;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24048;
    wire N__24045;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24037;
    wire N__24034;
    wire N__24031;
    wire N__24028;
    wire N__24025;
    wire N__24018;
    wire N__24015;
    wire N__24014;
    wire N__24013;
    wire N__24010;
    wire N__24005;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23993;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23976;
    wire N__23973;
    wire N__23972;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23957;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23945;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23928;
    wire N__23925;
    wire N__23924;
    wire N__23923;
    wire N__23920;
    wire N__23915;
    wire N__23910;
    wire N__23907;
    wire N__23906;
    wire N__23905;
    wire N__23902;
    wire N__23897;
    wire N__23892;
    wire N__23889;
    wire N__23888;
    wire N__23887;
    wire N__23884;
    wire N__23879;
    wire N__23874;
    wire N__23871;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23844;
    wire N__23841;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23814;
    wire N__23811;
    wire N__23810;
    wire N__23809;
    wire N__23806;
    wire N__23801;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23789;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23772;
    wire N__23769;
    wire N__23768;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23753;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23741;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23731;
    wire N__23724;
    wire N__23721;
    wire N__23720;
    wire N__23719;
    wire N__23716;
    wire N__23711;
    wire N__23706;
    wire N__23703;
    wire N__23702;
    wire N__23699;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23689;
    wire N__23682;
    wire N__23679;
    wire N__23678;
    wire N__23675;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23658;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23650;
    wire N__23645;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23633;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23616;
    wire N__23613;
    wire N__23612;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23597;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23585;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23568;
    wire N__23565;
    wire N__23564;
    wire N__23563;
    wire N__23560;
    wire N__23555;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23511;
    wire N__23510;
    wire N__23505;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23241;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23159;
    wire N__23158;
    wire N__23157;
    wire N__23156;
    wire N__23155;
    wire N__23154;
    wire N__23153;
    wire N__23152;
    wire N__23151;
    wire N__23150;
    wire N__23149;
    wire N__23148;
    wire N__23147;
    wire N__23146;
    wire N__23145;
    wire N__23128;
    wire N__23111;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23091;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23067;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23007;
    wire N__23004;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22832;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22816;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22791;
    wire N__22790;
    wire N__22787;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22773;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22752;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22714;
    wire N__22707;
    wire N__22706;
    wire N__22705;
    wire N__22704;
    wire N__22703;
    wire N__22702;
    wire N__22701;
    wire N__22700;
    wire N__22699;
    wire N__22698;
    wire N__22697;
    wire N__22696;
    wire N__22695;
    wire N__22694;
    wire N__22693;
    wire N__22692;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22668;
    wire N__22665;
    wire N__22664;
    wire N__22661;
    wire N__22660;
    wire N__22659;
    wire N__22658;
    wire N__22657;
    wire N__22656;
    wire N__22655;
    wire N__22654;
    wire N__22653;
    wire N__22652;
    wire N__22651;
    wire N__22650;
    wire N__22649;
    wire N__22648;
    wire N__22635;
    wire N__22632;
    wire N__22621;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22599;
    wire N__22596;
    wire N__22585;
    wire N__22582;
    wire N__22577;
    wire N__22574;
    wire N__22569;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22470;
    wire N__22467;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22437;
    wire N__22434;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22407;
    wire N__22404;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22392;
    wire N__22389;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22364;
    wire N__22361;
    wire N__22356;
    wire N__22353;
    wire N__22352;
    wire N__22347;
    wire N__22344;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22326;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22301;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22289;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22277;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22262;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22250;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22229;
    wire N__22228;
    wire N__22227;
    wire N__22226;
    wire N__22225;
    wire N__22224;
    wire N__22223;
    wire N__22222;
    wire N__22219;
    wire N__22218;
    wire N__22215;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22207;
    wire N__22204;
    wire N__22203;
    wire N__22200;
    wire N__22199;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22178;
    wire N__22161;
    wire N__22158;
    wire N__22157;
    wire N__22154;
    wire N__22149;
    wire N__22142;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22121;
    wire N__22118;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22076;
    wire N__22073;
    wire N__22072;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22045;
    wire N__22038;
    wire N__22035;
    wire N__22034;
    wire N__22031;
    wire N__22030;
    wire N__22027;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22003;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21986;
    wire N__21983;
    wire N__21982;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21924;
    wire N__21921;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21891;
    wire N__21888;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21860;
    wire N__21859;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21835;
    wire N__21828;
    wire N__21825;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21804;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21773;
    wire N__21770;
    wire N__21769;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21742;
    wire N__21735;
    wire N__21732;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21724;
    wire N__21721;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21687;
    wire N__21684;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21672;
    wire N__21669;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21654;
    wire N__21651;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21643;
    wire N__21640;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21622;
    wire N__21619;
    wire N__21612;
    wire N__21609;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21592;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21571;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21535;
    wire N__21530;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21477;
    wire N__21474;
    wire N__21469;
    wire N__21466;
    wire N__21459;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21437;
    wire N__21436;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21407;
    wire N__21402;
    wire N__21399;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21371;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21340;
    wire N__21337;
    wire N__21330;
    wire N__21327;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21312;
    wire N__21309;
    wire N__21308;
    wire N__21305;
    wire N__21302;
    wire N__21301;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21283;
    wire N__21278;
    wire N__21273;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21251;
    wire N__21248;
    wire N__21247;
    wire N__21244;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21220;
    wire N__21213;
    wire N__21210;
    wire N__21209;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21175;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21161;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21141;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21107;
    wire N__21106;
    wire N__21103;
    wire N__21098;
    wire N__21095;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21069;
    wire N__21066;
    wire N__21065;
    wire N__21064;
    wire N__21061;
    wire N__21056;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21035;
    wire N__21034;
    wire N__21031;
    wire N__21026;
    wire N__21023;
    wire N__21022;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21003;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20995;
    wire N__20994;
    wire N__20989;
    wire N__20984;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20957;
    wire N__20956;
    wire N__20953;
    wire N__20948;
    wire N__20943;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20931;
    wire N__20928;
    wire N__20927;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20900;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20882;
    wire N__20879;
    wire N__20878;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20862;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20844;
    wire N__20841;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20816;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20795;
    wire N__20792;
    wire N__20791;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20779;
    wire N__20776;
    wire N__20769;
    wire N__20766;
    wire N__20765;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20738;
    wire N__20733;
    wire N__20730;
    wire N__20729;
    wire N__20728;
    wire N__20727;
    wire N__20724;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20691;
    wire N__20688;
    wire N__20687;
    wire N__20684;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20663;
    wire N__20658;
    wire N__20655;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20647;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20591;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20567;
    wire N__20566;
    wire N__20565;
    wire N__20562;
    wire N__20561;
    wire N__20560;
    wire N__20559;
    wire N__20558;
    wire N__20557;
    wire N__20556;
    wire N__20555;
    wire N__20554;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20526;
    wire N__20525;
    wire N__20524;
    wire N__20523;
    wire N__20522;
    wire N__20521;
    wire N__20520;
    wire N__20519;
    wire N__20518;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20514;
    wire N__20513;
    wire N__20512;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20494;
    wire N__20483;
    wire N__20470;
    wire N__20467;
    wire N__20452;
    wire N__20441;
    wire N__20434;
    wire N__20431;
    wire N__20422;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20399;
    wire N__20398;
    wire N__20397;
    wire N__20396;
    wire N__20395;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20387;
    wire N__20386;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20378;
    wire N__20377;
    wire N__20376;
    wire N__20375;
    wire N__20374;
    wire N__20373;
    wire N__20372;
    wire N__20371;
    wire N__20370;
    wire N__20369;
    wire N__20368;
    wire N__20357;
    wire N__20356;
    wire N__20355;
    wire N__20354;
    wire N__20353;
    wire N__20352;
    wire N__20351;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20336;
    wire N__20333;
    wire N__20326;
    wire N__20317;
    wire N__20316;
    wire N__20315;
    wire N__20314;
    wire N__20311;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20287;
    wire N__20282;
    wire N__20277;
    wire N__20274;
    wire N__20269;
    wire N__20266;
    wire N__20255;
    wire N__20250;
    wire N__20245;
    wire N__20240;
    wire N__20229;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20214;
    wire N__20213;
    wire N__20210;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20195;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20166;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20105;
    wire N__20102;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20082;
    wire N__20079;
    wire N__20078;
    wire N__20075;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20055;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19964;
    wire N__19963;
    wire N__19962;
    wire N__19961;
    wire N__19960;
    wire N__19957;
    wire N__19948;
    wire N__19947;
    wire N__19946;
    wire N__19945;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19917;
    wire N__19914;
    wire N__19913;
    wire N__19908;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19875;
    wire N__19872;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19857;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19842;
    wire N__19839;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19824;
    wire N__19823;
    wire N__19822;
    wire N__19819;
    wire N__19814;
    wire N__19811;
    wire N__19806;
    wire N__19803;
    wire N__19802;
    wire N__19801;
    wire N__19798;
    wire N__19793;
    wire N__19790;
    wire N__19785;
    wire N__19784;
    wire N__19781;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19769;
    wire N__19766;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19754;
    wire N__19753;
    wire N__19750;
    wire N__19745;
    wire N__19742;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19703;
    wire N__19702;
    wire N__19701;
    wire N__19700;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19678;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19640;
    wire N__19639;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19363;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19344;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19332;
    wire N__19331;
    wire N__19330;
    wire N__19329;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19077;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19041;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire N__18996;
    wire N__18993;
    wire N__18990;
    wire N__18987;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18966;
    wire N__18963;
    wire N__18960;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18758;
    wire N__18757;
    wire N__18754;
    wire N__18753;
    wire N__18750;
    wire N__18741;
    wire N__18740;
    wire N__18739;
    wire N__18738;
    wire N__18737;
    wire N__18736;
    wire N__18735;
    wire N__18734;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18696;
    wire N__18687;
    wire N__18682;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18489;
    wire N__18486;
    wire N__18483;
    wire N__18480;
    wire N__18477;
    wire N__18474;
    wire N__18471;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18426;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire bfn_1_10_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire bfn_1_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire bfn_1_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire bfn_1_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire bfn_1_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire bfn_1_15_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ;
    wire \current_shift_inst.PI_CTRL.N_98_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_96_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire N_38_i_i;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_77_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.N_159 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire pwm_duty_input_7;
    wire pwm_duty_input_8;
    wire pwm_duty_input_6;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire pwm_duty_input_9;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire pwm_duty_input_4;
    wire pwm_duty_input_3;
    wire pwm_duty_input_5;
    wire rgb_drv_RNOZ0;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.N_46 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire bfn_3_17_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire bfn_3_18_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire bfn_3_19_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire bfn_3_20_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_5_15_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire bfn_5_16_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13_cascade_;
    wire bfn_7_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire bfn_7_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_7_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_7_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_7_26_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_7_27_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire bfn_7_28_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire il_max_comp1_c;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_8_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_8_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_8_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_8_14_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \current_shift_inst.control_input_18 ;
    wire bfn_8_15_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_8_16_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire s4_phy_c;
    wire GB_BUFFER_clock_output_0_THRU_CO;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire elapsed_time_ns_1_RNI68CN9_0_19_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire elapsed_time_ns_1_RNIK63T9_0_8_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire il_min_comp1_c;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.N_198_i ;
    wire \delay_measurement_inst.delay_hc_timer.N_199_i ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.N_1288_i ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire bfn_9_26_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire bfn_9_27_0_;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire bfn_9_28_0_;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire elapsed_time_ns_1_RNIU0DN9_0_20_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire elapsed_time_ns_1_RNIUVBN9_0_11_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12_cascade_;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.un1_start_g ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire bfn_10_26_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ;
    wire bfn_10_27_0_;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire bfn_10_28_0_;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire bfn_11_5_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_11_6_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_11_7_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_11_8_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_11_11_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_11_12_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire bfn_11_13_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire il_max_comp1_D1;
    wire il_min_comp1_D1;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire bfn_11_17_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire bfn_11_18_0_;
    wire \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_11_19_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire bfn_11_20_0_;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire s3_phy_c;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire bfn_11_24_0_;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire bfn_11_25_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire delay_hc_input_c_g;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_12_7_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_12_8_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire bfn_12_9_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_12_10_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_12_11_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_12_12_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_12_13_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire il_max_comp1_D2;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ;
    wire bfn_12_17_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire bfn_12_18_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_12_19_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_12_20_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire s1_phy_c;
    wire state_3;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ;
    wire \pll_inst.red_c_i ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire bfn_13_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire bfn_13_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_13_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_13_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire start_stop_c;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_162_i ;
    wire bfn_13_22_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_13_23_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.state_RNIE87FZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_13_24_0_;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_13_25_0_;
    wire \pwm_generator_inst.threshold_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire bfn_14_5_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_14_6_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_14_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_14_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_201_i ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21_cascade_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_14_11_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_14_12_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire bfn_14_13_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire bfn_14_18_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_14_19_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_14_20_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ;
    wire \pwm_generator_inst.N_16 ;
    wire N_19_1;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.threshold_0 ;
    wire state_ns_i_a3_1;
    wire T45_c;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.time_passed_RNIG7JF ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_200_i ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire elapsed_time_ns_1_RNIV8OBB_0_12_cascade_;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt20 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire elapsed_time_ns_1_RNI4EOBB_0_17_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire elapsed_time_ns_1_RNI3DOBB_0_16_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire bfn_15_13_0_;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_15_14_0_;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire bfn_15_15_0_;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_15_16_0_;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire \phase_controller_inst2.start_timer_tr_RNO_0_0 ;
    wire il_max_comp2_c;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire T12_c;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_16_8_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_16_9_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire bfn_16_10_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_16_11_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_16_12_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_16_13_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_16_14_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire T01_c;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire bfn_17_7_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_17_8_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_17_9_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_17_10_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire T23_c;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df30 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire bfn_17_15_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire bfn_17_16_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire bfn_17_17_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.N_162_i_g ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_17_19_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_17_20_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_17_21_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_17_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_163_i ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire elapsed_time_ns_1_RNI4FPBB_0_26_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire elapsed_time_ns_1_RNI5GPBB_0_27_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire elapsed_time_ns_1_RNI6HPBB_0_28_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire elapsed_time_ns_1_RNI3EPBB_0_25_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire elapsed_time_ns_1_RNI2DPBB_0_24_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_start_g ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire clock_output_0;
    wire red_c_g;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire _gnd_net_;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__24459),
            .RESETB(N__32172),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clock_output_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__35676),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__35581),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__23152,N__23160,N__23151,N__23158,N__23150,N__23157,N__23149,N__23159,N__23146,N__23153,N__23145,N__23154,N__23148,N__23155,N__23147,N__23156}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__35583,dangling_wire_45,N__35582}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__35664),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__35657),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__36015,N__36008,N__36013,N__36007,N__36014,N__36006,N__36016,N__36003,N__36009,N__36002,N__36010,N__36004,N__36011,N__36005,N__36012}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,N__35663,N__35660,dangling_wire_102,dangling_wire_103,dangling_wire_104,N__35658,N__35662,N__35659,N__35661}),
            .OHOLDTOP(),
            .O({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__35607),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__35591),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .ADDSUBBOT(),
            .A({dangling_wire_136,N__36017,N__36020,N__36018,N__36021,N__36019,N__19758,N__19806,N__19824,N__19785,N__20055,N__20105,N__20078,N__19842,N__19857,N__19875}),
            .C({dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}),
            .B({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,N__35597,N__35594,dangling_wire_160,dangling_wire_161,dangling_wire_162,N__35592,N__35596,N__35593,N__35595}),
            .OHOLDTOP(),
            .O({dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__35671),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__35668),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .ADDSUBBOT(),
            .A({dangling_wire_185,N__23110,N__22875,N__22899,N__22926,N__22953,N__23067,N__22977,N__23004,N__23031,N__22434,N__22466,N__22494,N__22518,N__22539,N__24387}),
            .C({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .B({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__35670,dangling_wire_215,N__35669}),
            .OHOLDTOP(),
            .O({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__48637),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__48639),
            .DIN(N__48638),
            .DOUT(N__48637),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__48639),
            .PADOUT(N__48638),
            .PADIN(N__48637),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clock_output_obuf_iopad (
            .OE(N__48628),
            .DIN(N__48627),
            .DOUT(N__48626),
            .PACKAGEPIN(clock_output));
    defparam clock_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam clock_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO clock_output_obuf_preio (
            .PADOEN(N__48628),
            .PADOUT(N__48627),
            .PADIN(N__48626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24477),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__48619),
            .DIN(N__48618),
            .DOUT(N__48617),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__48619),
            .PADOUT(N__48618),
            .PADIN(N__48617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__39537),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__48610),
            .DIN(N__48609),
            .DOUT(N__48608),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__48610),
            .PADOUT(N__48609),
            .PADIN(N__48608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__48601),
            .DIN(N__48600),
            .DOUT(N__48599),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__48601),
            .PADOUT(N__48600),
            .PADIN(N__48599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__48592),
            .DIN(N__48591),
            .DOUT(N__48590),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__48592),
            .PADOUT(N__48591),
            .PADIN(N__48590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__41892),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__48583),
            .DIN(N__48582),
            .DOUT(N__48581),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__48583),
            .PADOUT(N__48582),
            .PADIN(N__48581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33489),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__48574),
            .DIN(N__48573),
            .DOUT(N__48572),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__48574),
            .PADOUT(N__48573),
            .PADIN(N__48572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__48565),
            .DIN(N__48564),
            .DOUT(N__48563),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__48565),
            .PADOUT(N__48564),
            .PADIN(N__48563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33426),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__48556),
            .DIN(N__48555),
            .DOUT(N__48554),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__48556),
            .PADOUT(N__48555),
            .PADIN(N__48554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__38433),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__48547),
            .DIN(N__48546),
            .DOUT(N__48545),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__48547),
            .PADOUT(N__48546),
            .PADIN(N__48545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__48538),
            .DIN(N__48537),
            .DOUT(N__48536),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__48538),
            .PADOUT(N__48537),
            .PADIN(N__48536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31797),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__48529),
            .DIN(N__48528),
            .DOUT(N__48527),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__48529),
            .PADOUT(N__48528),
            .PADIN(N__48527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24360),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__48520),
            .DIN(N__48519),
            .DOUT(N__48518),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__48520),
            .PADOUT(N__48519),
            .PADIN(N__48518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__48511),
            .DIN(N__48510),
            .DOUT(N__48509),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__48511),
            .PADOUT(N__48510),
            .PADIN(N__48509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29403),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__48502),
            .DIN(N__48501),
            .DOUT(N__48500),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__48502),
            .PADOUT(N__48501),
            .PADIN(N__48500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35769),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__48493),
            .DIN(N__48492),
            .DOUT(N__48491),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__48493),
            .PADOUT(N__48492),
            .PADIN(N__48491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__48484),
            .DIN(N__48483),
            .DOUT(N__48482),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__48484),
            .PADOUT(N__48483),
            .PADIN(N__48482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11559 (
            .O(N__48465),
            .I(N__48460));
    InMux I__11558 (
            .O(N__48464),
            .I(N__48457));
    InMux I__11557 (
            .O(N__48463),
            .I(N__48454));
    LocalMux I__11556 (
            .O(N__48460),
            .I(N__48449));
    LocalMux I__11555 (
            .O(N__48457),
            .I(N__48449));
    LocalMux I__11554 (
            .O(N__48454),
            .I(N__48445));
    Span4Mux_v I__11553 (
            .O(N__48449),
            .I(N__48442));
    InMux I__11552 (
            .O(N__48448),
            .I(N__48439));
    Span4Mux_v I__11551 (
            .O(N__48445),
            .I(N__48436));
    Sp12to4 I__11550 (
            .O(N__48442),
            .I(N__48431));
    LocalMux I__11549 (
            .O(N__48439),
            .I(N__48431));
    Odrv4 I__11548 (
            .O(N__48436),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv12 I__11547 (
            .O(N__48431),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__11546 (
            .O(N__48426),
            .I(N__48422));
    InMux I__11545 (
            .O(N__48425),
            .I(N__48418));
    LocalMux I__11544 (
            .O(N__48422),
            .I(N__48415));
    InMux I__11543 (
            .O(N__48421),
            .I(N__48412));
    LocalMux I__11542 (
            .O(N__48418),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    Odrv12 I__11541 (
            .O(N__48415),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    LocalMux I__11540 (
            .O(N__48412),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__11539 (
            .O(N__48405),
            .I(N__48402));
    LocalMux I__11538 (
            .O(N__48402),
            .I(N__48397));
    InMux I__11537 (
            .O(N__48401),
            .I(N__48394));
    InMux I__11536 (
            .O(N__48400),
            .I(N__48391));
    Span4Mux_v I__11535 (
            .O(N__48397),
            .I(N__48388));
    LocalMux I__11534 (
            .O(N__48394),
            .I(N__48385));
    LocalMux I__11533 (
            .O(N__48391),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv4 I__11532 (
            .O(N__48388),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv4 I__11531 (
            .O(N__48385),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    InMux I__11530 (
            .O(N__48378),
            .I(N__48373));
    InMux I__11529 (
            .O(N__48377),
            .I(N__48370));
    InMux I__11528 (
            .O(N__48376),
            .I(N__48367));
    LocalMux I__11527 (
            .O(N__48373),
            .I(N__48362));
    LocalMux I__11526 (
            .O(N__48370),
            .I(N__48362));
    LocalMux I__11525 (
            .O(N__48367),
            .I(N__48359));
    Span12Mux_h I__11524 (
            .O(N__48362),
            .I(N__48355));
    Span4Mux_h I__11523 (
            .O(N__48359),
            .I(N__48352));
    InMux I__11522 (
            .O(N__48358),
            .I(N__48349));
    Odrv12 I__11521 (
            .O(N__48355),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__11520 (
            .O(N__48352),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    LocalMux I__11519 (
            .O(N__48349),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__11518 (
            .O(N__48342),
            .I(N__48315));
    InMux I__11517 (
            .O(N__48341),
            .I(N__48315));
    InMux I__11516 (
            .O(N__48340),
            .I(N__48315));
    CascadeMux I__11515 (
            .O(N__48339),
            .I(N__48311));
    InMux I__11514 (
            .O(N__48338),
            .I(N__48302));
    InMux I__11513 (
            .O(N__48337),
            .I(N__48279));
    InMux I__11512 (
            .O(N__48336),
            .I(N__48279));
    InMux I__11511 (
            .O(N__48335),
            .I(N__48272));
    InMux I__11510 (
            .O(N__48334),
            .I(N__48272));
    InMux I__11509 (
            .O(N__48333),
            .I(N__48272));
    InMux I__11508 (
            .O(N__48332),
            .I(N__48269));
    InMux I__11507 (
            .O(N__48331),
            .I(N__48234));
    InMux I__11506 (
            .O(N__48330),
            .I(N__48234));
    InMux I__11505 (
            .O(N__48329),
            .I(N__48234));
    InMux I__11504 (
            .O(N__48328),
            .I(N__48234));
    InMux I__11503 (
            .O(N__48327),
            .I(N__48234));
    InMux I__11502 (
            .O(N__48326),
            .I(N__48234));
    InMux I__11501 (
            .O(N__48325),
            .I(N__48231));
    InMux I__11500 (
            .O(N__48324),
            .I(N__48220));
    InMux I__11499 (
            .O(N__48323),
            .I(N__48220));
    InMux I__11498 (
            .O(N__48322),
            .I(N__48217));
    LocalMux I__11497 (
            .O(N__48315),
            .I(N__48214));
    InMux I__11496 (
            .O(N__48314),
            .I(N__48201));
    InMux I__11495 (
            .O(N__48311),
            .I(N__48201));
    InMux I__11494 (
            .O(N__48310),
            .I(N__48201));
    InMux I__11493 (
            .O(N__48309),
            .I(N__48201));
    InMux I__11492 (
            .O(N__48308),
            .I(N__48201));
    InMux I__11491 (
            .O(N__48307),
            .I(N__48201));
    InMux I__11490 (
            .O(N__48306),
            .I(N__48196));
    InMux I__11489 (
            .O(N__48305),
            .I(N__48196));
    LocalMux I__11488 (
            .O(N__48302),
            .I(N__48193));
    InMux I__11487 (
            .O(N__48301),
            .I(N__48173));
    InMux I__11486 (
            .O(N__48300),
            .I(N__48173));
    InMux I__11485 (
            .O(N__48299),
            .I(N__48173));
    InMux I__11484 (
            .O(N__48298),
            .I(N__48173));
    InMux I__11483 (
            .O(N__48297),
            .I(N__48173));
    InMux I__11482 (
            .O(N__48296),
            .I(N__48166));
    InMux I__11481 (
            .O(N__48295),
            .I(N__48166));
    InMux I__11480 (
            .O(N__48294),
            .I(N__48166));
    InMux I__11479 (
            .O(N__48293),
            .I(N__48163));
    InMux I__11478 (
            .O(N__48292),
            .I(N__48152));
    InMux I__11477 (
            .O(N__48291),
            .I(N__48152));
    InMux I__11476 (
            .O(N__48290),
            .I(N__48152));
    InMux I__11475 (
            .O(N__48289),
            .I(N__48152));
    InMux I__11474 (
            .O(N__48288),
            .I(N__48152));
    InMux I__11473 (
            .O(N__48287),
            .I(N__48143));
    InMux I__11472 (
            .O(N__48286),
            .I(N__48143));
    InMux I__11471 (
            .O(N__48285),
            .I(N__48143));
    InMux I__11470 (
            .O(N__48284),
            .I(N__48143));
    LocalMux I__11469 (
            .O(N__48279),
            .I(N__48138));
    LocalMux I__11468 (
            .O(N__48272),
            .I(N__48138));
    LocalMux I__11467 (
            .O(N__48269),
            .I(N__48135));
    InMux I__11466 (
            .O(N__48268),
            .I(N__48132));
    InMux I__11465 (
            .O(N__48267),
            .I(N__48121));
    InMux I__11464 (
            .O(N__48266),
            .I(N__48121));
    InMux I__11463 (
            .O(N__48265),
            .I(N__48121));
    InMux I__11462 (
            .O(N__48264),
            .I(N__48121));
    InMux I__11461 (
            .O(N__48263),
            .I(N__48121));
    InMux I__11460 (
            .O(N__48262),
            .I(N__48115));
    InMux I__11459 (
            .O(N__48261),
            .I(N__48106));
    InMux I__11458 (
            .O(N__48260),
            .I(N__48106));
    InMux I__11457 (
            .O(N__48259),
            .I(N__48106));
    InMux I__11456 (
            .O(N__48258),
            .I(N__48106));
    InMux I__11455 (
            .O(N__48257),
            .I(N__48101));
    InMux I__11454 (
            .O(N__48256),
            .I(N__48101));
    InMux I__11453 (
            .O(N__48255),
            .I(N__48092));
    InMux I__11452 (
            .O(N__48254),
            .I(N__48092));
    InMux I__11451 (
            .O(N__48253),
            .I(N__48092));
    InMux I__11450 (
            .O(N__48252),
            .I(N__48092));
    InMux I__11449 (
            .O(N__48251),
            .I(N__48081));
    InMux I__11448 (
            .O(N__48250),
            .I(N__48081));
    InMux I__11447 (
            .O(N__48249),
            .I(N__48081));
    InMux I__11446 (
            .O(N__48248),
            .I(N__48081));
    InMux I__11445 (
            .O(N__48247),
            .I(N__48081));
    LocalMux I__11444 (
            .O(N__48234),
            .I(N__48078));
    LocalMux I__11443 (
            .O(N__48231),
            .I(N__48075));
    InMux I__11442 (
            .O(N__48230),
            .I(N__48060));
    InMux I__11441 (
            .O(N__48229),
            .I(N__48060));
    InMux I__11440 (
            .O(N__48228),
            .I(N__48060));
    InMux I__11439 (
            .O(N__48227),
            .I(N__48060));
    InMux I__11438 (
            .O(N__48226),
            .I(N__48060));
    InMux I__11437 (
            .O(N__48225),
            .I(N__48060));
    LocalMux I__11436 (
            .O(N__48220),
            .I(N__48057));
    LocalMux I__11435 (
            .O(N__48217),
            .I(N__48050));
    Span4Mux_h I__11434 (
            .O(N__48214),
            .I(N__48050));
    LocalMux I__11433 (
            .O(N__48201),
            .I(N__48050));
    LocalMux I__11432 (
            .O(N__48196),
            .I(N__48045));
    Span4Mux_v I__11431 (
            .O(N__48193),
            .I(N__48045));
    InMux I__11430 (
            .O(N__48192),
            .I(N__48034));
    InMux I__11429 (
            .O(N__48191),
            .I(N__48034));
    InMux I__11428 (
            .O(N__48190),
            .I(N__48034));
    InMux I__11427 (
            .O(N__48189),
            .I(N__48031));
    InMux I__11426 (
            .O(N__48188),
            .I(N__48026));
    InMux I__11425 (
            .O(N__48187),
            .I(N__48026));
    InMux I__11424 (
            .O(N__48186),
            .I(N__48019));
    InMux I__11423 (
            .O(N__48185),
            .I(N__48019));
    InMux I__11422 (
            .O(N__48184),
            .I(N__48019));
    LocalMux I__11421 (
            .O(N__48173),
            .I(N__48014));
    LocalMux I__11420 (
            .O(N__48166),
            .I(N__48014));
    LocalMux I__11419 (
            .O(N__48163),
            .I(N__48011));
    LocalMux I__11418 (
            .O(N__48152),
            .I(N__48004));
    LocalMux I__11417 (
            .O(N__48143),
            .I(N__48004));
    Span4Mux_v I__11416 (
            .O(N__48138),
            .I(N__48004));
    Span4Mux_h I__11415 (
            .O(N__48135),
            .I(N__47999));
    LocalMux I__11414 (
            .O(N__48132),
            .I(N__47999));
    LocalMux I__11413 (
            .O(N__48121),
            .I(N__47996));
    InMux I__11412 (
            .O(N__48120),
            .I(N__47993));
    InMux I__11411 (
            .O(N__48119),
            .I(N__47988));
    InMux I__11410 (
            .O(N__48118),
            .I(N__47988));
    LocalMux I__11409 (
            .O(N__48115),
            .I(N__47985));
    LocalMux I__11408 (
            .O(N__48106),
            .I(N__47978));
    LocalMux I__11407 (
            .O(N__48101),
            .I(N__47978));
    LocalMux I__11406 (
            .O(N__48092),
            .I(N__47978));
    LocalMux I__11405 (
            .O(N__48081),
            .I(N__47971));
    Span4Mux_v I__11404 (
            .O(N__48078),
            .I(N__47971));
    Span4Mux_v I__11403 (
            .O(N__48075),
            .I(N__47971));
    InMux I__11402 (
            .O(N__48074),
            .I(N__47966));
    InMux I__11401 (
            .O(N__48073),
            .I(N__47966));
    LocalMux I__11400 (
            .O(N__48060),
            .I(N__47957));
    Span4Mux_v I__11399 (
            .O(N__48057),
            .I(N__47957));
    Span4Mux_v I__11398 (
            .O(N__48050),
            .I(N__47957));
    Span4Mux_v I__11397 (
            .O(N__48045),
            .I(N__47957));
    InMux I__11396 (
            .O(N__48044),
            .I(N__47954));
    InMux I__11395 (
            .O(N__48043),
            .I(N__47947));
    InMux I__11394 (
            .O(N__48042),
            .I(N__47947));
    InMux I__11393 (
            .O(N__48041),
            .I(N__47947));
    LocalMux I__11392 (
            .O(N__48034),
            .I(N__47944));
    LocalMux I__11391 (
            .O(N__48031),
            .I(N__47939));
    LocalMux I__11390 (
            .O(N__48026),
            .I(N__47939));
    LocalMux I__11389 (
            .O(N__48019),
            .I(N__47928));
    Span4Mux_v I__11388 (
            .O(N__48014),
            .I(N__47928));
    Span4Mux_h I__11387 (
            .O(N__48011),
            .I(N__47928));
    Span4Mux_h I__11386 (
            .O(N__48004),
            .I(N__47928));
    Span4Mux_h I__11385 (
            .O(N__47999),
            .I(N__47928));
    Span12Mux_h I__11384 (
            .O(N__47996),
            .I(N__47925));
    LocalMux I__11383 (
            .O(N__47993),
            .I(N__47914));
    LocalMux I__11382 (
            .O(N__47988),
            .I(N__47914));
    Span4Mux_h I__11381 (
            .O(N__47985),
            .I(N__47914));
    Span4Mux_v I__11380 (
            .O(N__47978),
            .I(N__47914));
    Span4Mux_h I__11379 (
            .O(N__47971),
            .I(N__47914));
    LocalMux I__11378 (
            .O(N__47966),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11377 (
            .O(N__47957),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11376 (
            .O(N__47954),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11375 (
            .O(N__47947),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11374 (
            .O(N__47944),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11373 (
            .O(N__47939),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11372 (
            .O(N__47928),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__11371 (
            .O(N__47925),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11370 (
            .O(N__47914),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    CascadeMux I__11369 (
            .O(N__47895),
            .I(N__47892));
    InMux I__11368 (
            .O(N__47892),
            .I(N__47886));
    InMux I__11367 (
            .O(N__47891),
            .I(N__47886));
    LocalMux I__11366 (
            .O(N__47886),
            .I(N__47883));
    Span4Mux_h I__11365 (
            .O(N__47883),
            .I(N__47880));
    Odrv4 I__11364 (
            .O(N__47880),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ));
    CEMux I__11363 (
            .O(N__47877),
            .I(N__47870));
    CEMux I__11362 (
            .O(N__47876),
            .I(N__47866));
    CEMux I__11361 (
            .O(N__47875),
            .I(N__47863));
    InMux I__11360 (
            .O(N__47874),
            .I(N__47858));
    CEMux I__11359 (
            .O(N__47873),
            .I(N__47855));
    LocalMux I__11358 (
            .O(N__47870),
            .I(N__47852));
    CEMux I__11357 (
            .O(N__47869),
            .I(N__47844));
    LocalMux I__11356 (
            .O(N__47866),
            .I(N__47816));
    LocalMux I__11355 (
            .O(N__47863),
            .I(N__47812));
    CEMux I__11354 (
            .O(N__47862),
            .I(N__47808));
    CEMux I__11353 (
            .O(N__47861),
            .I(N__47805));
    LocalMux I__11352 (
            .O(N__47858),
            .I(N__47802));
    LocalMux I__11351 (
            .O(N__47855),
            .I(N__47799));
    Span4Mux_h I__11350 (
            .O(N__47852),
            .I(N__47796));
    CEMux I__11349 (
            .O(N__47851),
            .I(N__47793));
    InMux I__11348 (
            .O(N__47850),
            .I(N__47784));
    InMux I__11347 (
            .O(N__47849),
            .I(N__47784));
    InMux I__11346 (
            .O(N__47848),
            .I(N__47784));
    InMux I__11345 (
            .O(N__47847),
            .I(N__47784));
    LocalMux I__11344 (
            .O(N__47844),
            .I(N__47781));
    InMux I__11343 (
            .O(N__47843),
            .I(N__47770));
    InMux I__11342 (
            .O(N__47842),
            .I(N__47770));
    InMux I__11341 (
            .O(N__47841),
            .I(N__47770));
    InMux I__11340 (
            .O(N__47840),
            .I(N__47761));
    InMux I__11339 (
            .O(N__47839),
            .I(N__47761));
    InMux I__11338 (
            .O(N__47838),
            .I(N__47761));
    InMux I__11337 (
            .O(N__47837),
            .I(N__47761));
    InMux I__11336 (
            .O(N__47836),
            .I(N__47752));
    InMux I__11335 (
            .O(N__47835),
            .I(N__47752));
    InMux I__11334 (
            .O(N__47834),
            .I(N__47752));
    InMux I__11333 (
            .O(N__47833),
            .I(N__47752));
    InMux I__11332 (
            .O(N__47832),
            .I(N__47743));
    InMux I__11331 (
            .O(N__47831),
            .I(N__47743));
    InMux I__11330 (
            .O(N__47830),
            .I(N__47743));
    InMux I__11329 (
            .O(N__47829),
            .I(N__47743));
    InMux I__11328 (
            .O(N__47828),
            .I(N__47736));
    InMux I__11327 (
            .O(N__47827),
            .I(N__47736));
    InMux I__11326 (
            .O(N__47826),
            .I(N__47736));
    CEMux I__11325 (
            .O(N__47825),
            .I(N__47732));
    CEMux I__11324 (
            .O(N__47824),
            .I(N__47729));
    CEMux I__11323 (
            .O(N__47823),
            .I(N__47726));
    InMux I__11322 (
            .O(N__47822),
            .I(N__47717));
    InMux I__11321 (
            .O(N__47821),
            .I(N__47717));
    InMux I__11320 (
            .O(N__47820),
            .I(N__47717));
    InMux I__11319 (
            .O(N__47819),
            .I(N__47717));
    Span4Mux_v I__11318 (
            .O(N__47816),
            .I(N__47714));
    CEMux I__11317 (
            .O(N__47815),
            .I(N__47711));
    Span4Mux_v I__11316 (
            .O(N__47812),
            .I(N__47708));
    CEMux I__11315 (
            .O(N__47811),
            .I(N__47705));
    LocalMux I__11314 (
            .O(N__47808),
            .I(N__47702));
    LocalMux I__11313 (
            .O(N__47805),
            .I(N__47699));
    Span4Mux_v I__11312 (
            .O(N__47802),
            .I(N__47696));
    Span4Mux_h I__11311 (
            .O(N__47799),
            .I(N__47685));
    Span4Mux_h I__11310 (
            .O(N__47796),
            .I(N__47685));
    LocalMux I__11309 (
            .O(N__47793),
            .I(N__47685));
    LocalMux I__11308 (
            .O(N__47784),
            .I(N__47685));
    Span4Mux_v I__11307 (
            .O(N__47781),
            .I(N__47685));
    InMux I__11306 (
            .O(N__47780),
            .I(N__47676));
    InMux I__11305 (
            .O(N__47779),
            .I(N__47676));
    InMux I__11304 (
            .O(N__47778),
            .I(N__47676));
    InMux I__11303 (
            .O(N__47777),
            .I(N__47676));
    LocalMux I__11302 (
            .O(N__47770),
            .I(N__47671));
    LocalMux I__11301 (
            .O(N__47761),
            .I(N__47671));
    LocalMux I__11300 (
            .O(N__47752),
            .I(N__47664));
    LocalMux I__11299 (
            .O(N__47743),
            .I(N__47664));
    LocalMux I__11298 (
            .O(N__47736),
            .I(N__47664));
    CEMux I__11297 (
            .O(N__47735),
            .I(N__47661));
    LocalMux I__11296 (
            .O(N__47732),
            .I(N__47656));
    LocalMux I__11295 (
            .O(N__47729),
            .I(N__47656));
    LocalMux I__11294 (
            .O(N__47726),
            .I(N__47653));
    LocalMux I__11293 (
            .O(N__47717),
            .I(N__47648));
    Span4Mux_h I__11292 (
            .O(N__47714),
            .I(N__47648));
    LocalMux I__11291 (
            .O(N__47711),
            .I(N__47645));
    Span4Mux_h I__11290 (
            .O(N__47708),
            .I(N__47640));
    LocalMux I__11289 (
            .O(N__47705),
            .I(N__47640));
    Span4Mux_v I__11288 (
            .O(N__47702),
            .I(N__47635));
    Span4Mux_h I__11287 (
            .O(N__47699),
            .I(N__47635));
    Span4Mux_h I__11286 (
            .O(N__47696),
            .I(N__47632));
    Span4Mux_v I__11285 (
            .O(N__47685),
            .I(N__47623));
    LocalMux I__11284 (
            .O(N__47676),
            .I(N__47623));
    Span4Mux_v I__11283 (
            .O(N__47671),
            .I(N__47623));
    Span4Mux_v I__11282 (
            .O(N__47664),
            .I(N__47623));
    LocalMux I__11281 (
            .O(N__47661),
            .I(N__47618));
    Span12Mux_h I__11280 (
            .O(N__47656),
            .I(N__47618));
    Span4Mux_v I__11279 (
            .O(N__47653),
            .I(N__47613));
    Span4Mux_h I__11278 (
            .O(N__47648),
            .I(N__47613));
    Span4Mux_h I__11277 (
            .O(N__47645),
            .I(N__47610));
    Sp12to4 I__11276 (
            .O(N__47640),
            .I(N__47607));
    Span4Mux_h I__11275 (
            .O(N__47635),
            .I(N__47604));
    Span4Mux_h I__11274 (
            .O(N__47632),
            .I(N__47601));
    Span4Mux_h I__11273 (
            .O(N__47623),
            .I(N__47598));
    Odrv12 I__11272 (
            .O(N__47618),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11271 (
            .O(N__47613),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11270 (
            .O(N__47610),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv12 I__11269 (
            .O(N__47607),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11268 (
            .O(N__47604),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11267 (
            .O(N__47601),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11266 (
            .O(N__47598),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__11265 (
            .O(N__47583),
            .I(N__47580));
    LocalMux I__11264 (
            .O(N__47580),
            .I(N__47577));
    Span4Mux_v I__11263 (
            .O(N__47577),
            .I(N__47573));
    InMux I__11262 (
            .O(N__47576),
            .I(N__47570));
    Span4Mux_h I__11261 (
            .O(N__47573),
            .I(N__47567));
    LocalMux I__11260 (
            .O(N__47570),
            .I(N__47564));
    Odrv4 I__11259 (
            .O(N__47567),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__11258 (
            .O(N__47564),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__11257 (
            .O(N__47559),
            .I(N__47556));
    LocalMux I__11256 (
            .O(N__47556),
            .I(N__47413));
    ClkMux I__11255 (
            .O(N__47555),
            .I(N__47127));
    ClkMux I__11254 (
            .O(N__47554),
            .I(N__47127));
    ClkMux I__11253 (
            .O(N__47553),
            .I(N__47127));
    ClkMux I__11252 (
            .O(N__47552),
            .I(N__47127));
    ClkMux I__11251 (
            .O(N__47551),
            .I(N__47127));
    ClkMux I__11250 (
            .O(N__47550),
            .I(N__47127));
    ClkMux I__11249 (
            .O(N__47549),
            .I(N__47127));
    ClkMux I__11248 (
            .O(N__47548),
            .I(N__47127));
    ClkMux I__11247 (
            .O(N__47547),
            .I(N__47127));
    ClkMux I__11246 (
            .O(N__47546),
            .I(N__47127));
    ClkMux I__11245 (
            .O(N__47545),
            .I(N__47127));
    ClkMux I__11244 (
            .O(N__47544),
            .I(N__47127));
    ClkMux I__11243 (
            .O(N__47543),
            .I(N__47127));
    ClkMux I__11242 (
            .O(N__47542),
            .I(N__47127));
    ClkMux I__11241 (
            .O(N__47541),
            .I(N__47127));
    ClkMux I__11240 (
            .O(N__47540),
            .I(N__47127));
    ClkMux I__11239 (
            .O(N__47539),
            .I(N__47127));
    ClkMux I__11238 (
            .O(N__47538),
            .I(N__47127));
    ClkMux I__11237 (
            .O(N__47537),
            .I(N__47127));
    ClkMux I__11236 (
            .O(N__47536),
            .I(N__47127));
    ClkMux I__11235 (
            .O(N__47535),
            .I(N__47127));
    ClkMux I__11234 (
            .O(N__47534),
            .I(N__47127));
    ClkMux I__11233 (
            .O(N__47533),
            .I(N__47127));
    ClkMux I__11232 (
            .O(N__47532),
            .I(N__47127));
    ClkMux I__11231 (
            .O(N__47531),
            .I(N__47127));
    ClkMux I__11230 (
            .O(N__47530),
            .I(N__47127));
    ClkMux I__11229 (
            .O(N__47529),
            .I(N__47127));
    ClkMux I__11228 (
            .O(N__47528),
            .I(N__47127));
    ClkMux I__11227 (
            .O(N__47527),
            .I(N__47127));
    ClkMux I__11226 (
            .O(N__47526),
            .I(N__47127));
    ClkMux I__11225 (
            .O(N__47525),
            .I(N__47127));
    ClkMux I__11224 (
            .O(N__47524),
            .I(N__47127));
    ClkMux I__11223 (
            .O(N__47523),
            .I(N__47127));
    ClkMux I__11222 (
            .O(N__47522),
            .I(N__47127));
    ClkMux I__11221 (
            .O(N__47521),
            .I(N__47127));
    ClkMux I__11220 (
            .O(N__47520),
            .I(N__47127));
    ClkMux I__11219 (
            .O(N__47519),
            .I(N__47127));
    ClkMux I__11218 (
            .O(N__47518),
            .I(N__47127));
    ClkMux I__11217 (
            .O(N__47517),
            .I(N__47127));
    ClkMux I__11216 (
            .O(N__47516),
            .I(N__47127));
    ClkMux I__11215 (
            .O(N__47515),
            .I(N__47127));
    ClkMux I__11214 (
            .O(N__47514),
            .I(N__47127));
    ClkMux I__11213 (
            .O(N__47513),
            .I(N__47127));
    ClkMux I__11212 (
            .O(N__47512),
            .I(N__47127));
    ClkMux I__11211 (
            .O(N__47511),
            .I(N__47127));
    ClkMux I__11210 (
            .O(N__47510),
            .I(N__47127));
    ClkMux I__11209 (
            .O(N__47509),
            .I(N__47127));
    ClkMux I__11208 (
            .O(N__47508),
            .I(N__47127));
    ClkMux I__11207 (
            .O(N__47507),
            .I(N__47127));
    ClkMux I__11206 (
            .O(N__47506),
            .I(N__47127));
    ClkMux I__11205 (
            .O(N__47505),
            .I(N__47127));
    ClkMux I__11204 (
            .O(N__47504),
            .I(N__47127));
    ClkMux I__11203 (
            .O(N__47503),
            .I(N__47127));
    ClkMux I__11202 (
            .O(N__47502),
            .I(N__47127));
    ClkMux I__11201 (
            .O(N__47501),
            .I(N__47127));
    ClkMux I__11200 (
            .O(N__47500),
            .I(N__47127));
    ClkMux I__11199 (
            .O(N__47499),
            .I(N__47127));
    ClkMux I__11198 (
            .O(N__47498),
            .I(N__47127));
    ClkMux I__11197 (
            .O(N__47497),
            .I(N__47127));
    ClkMux I__11196 (
            .O(N__47496),
            .I(N__47127));
    ClkMux I__11195 (
            .O(N__47495),
            .I(N__47127));
    ClkMux I__11194 (
            .O(N__47494),
            .I(N__47127));
    ClkMux I__11193 (
            .O(N__47493),
            .I(N__47127));
    ClkMux I__11192 (
            .O(N__47492),
            .I(N__47127));
    ClkMux I__11191 (
            .O(N__47491),
            .I(N__47127));
    ClkMux I__11190 (
            .O(N__47490),
            .I(N__47127));
    ClkMux I__11189 (
            .O(N__47489),
            .I(N__47127));
    ClkMux I__11188 (
            .O(N__47488),
            .I(N__47127));
    ClkMux I__11187 (
            .O(N__47487),
            .I(N__47127));
    ClkMux I__11186 (
            .O(N__47486),
            .I(N__47127));
    ClkMux I__11185 (
            .O(N__47485),
            .I(N__47127));
    ClkMux I__11184 (
            .O(N__47484),
            .I(N__47127));
    ClkMux I__11183 (
            .O(N__47483),
            .I(N__47127));
    ClkMux I__11182 (
            .O(N__47482),
            .I(N__47127));
    ClkMux I__11181 (
            .O(N__47481),
            .I(N__47127));
    ClkMux I__11180 (
            .O(N__47480),
            .I(N__47127));
    ClkMux I__11179 (
            .O(N__47479),
            .I(N__47127));
    ClkMux I__11178 (
            .O(N__47478),
            .I(N__47127));
    ClkMux I__11177 (
            .O(N__47477),
            .I(N__47127));
    ClkMux I__11176 (
            .O(N__47476),
            .I(N__47127));
    ClkMux I__11175 (
            .O(N__47475),
            .I(N__47127));
    ClkMux I__11174 (
            .O(N__47474),
            .I(N__47127));
    ClkMux I__11173 (
            .O(N__47473),
            .I(N__47127));
    ClkMux I__11172 (
            .O(N__47472),
            .I(N__47127));
    ClkMux I__11171 (
            .O(N__47471),
            .I(N__47127));
    ClkMux I__11170 (
            .O(N__47470),
            .I(N__47127));
    ClkMux I__11169 (
            .O(N__47469),
            .I(N__47127));
    ClkMux I__11168 (
            .O(N__47468),
            .I(N__47127));
    ClkMux I__11167 (
            .O(N__47467),
            .I(N__47127));
    ClkMux I__11166 (
            .O(N__47466),
            .I(N__47127));
    ClkMux I__11165 (
            .O(N__47465),
            .I(N__47127));
    ClkMux I__11164 (
            .O(N__47464),
            .I(N__47127));
    ClkMux I__11163 (
            .O(N__47463),
            .I(N__47127));
    ClkMux I__11162 (
            .O(N__47462),
            .I(N__47127));
    ClkMux I__11161 (
            .O(N__47461),
            .I(N__47127));
    ClkMux I__11160 (
            .O(N__47460),
            .I(N__47127));
    ClkMux I__11159 (
            .O(N__47459),
            .I(N__47127));
    ClkMux I__11158 (
            .O(N__47458),
            .I(N__47127));
    ClkMux I__11157 (
            .O(N__47457),
            .I(N__47127));
    ClkMux I__11156 (
            .O(N__47456),
            .I(N__47127));
    ClkMux I__11155 (
            .O(N__47455),
            .I(N__47127));
    ClkMux I__11154 (
            .O(N__47454),
            .I(N__47127));
    ClkMux I__11153 (
            .O(N__47453),
            .I(N__47127));
    ClkMux I__11152 (
            .O(N__47452),
            .I(N__47127));
    ClkMux I__11151 (
            .O(N__47451),
            .I(N__47127));
    ClkMux I__11150 (
            .O(N__47450),
            .I(N__47127));
    ClkMux I__11149 (
            .O(N__47449),
            .I(N__47127));
    ClkMux I__11148 (
            .O(N__47448),
            .I(N__47127));
    ClkMux I__11147 (
            .O(N__47447),
            .I(N__47127));
    ClkMux I__11146 (
            .O(N__47446),
            .I(N__47127));
    ClkMux I__11145 (
            .O(N__47445),
            .I(N__47127));
    ClkMux I__11144 (
            .O(N__47444),
            .I(N__47127));
    ClkMux I__11143 (
            .O(N__47443),
            .I(N__47127));
    ClkMux I__11142 (
            .O(N__47442),
            .I(N__47127));
    ClkMux I__11141 (
            .O(N__47441),
            .I(N__47127));
    ClkMux I__11140 (
            .O(N__47440),
            .I(N__47127));
    ClkMux I__11139 (
            .O(N__47439),
            .I(N__47127));
    ClkMux I__11138 (
            .O(N__47438),
            .I(N__47127));
    ClkMux I__11137 (
            .O(N__47437),
            .I(N__47127));
    ClkMux I__11136 (
            .O(N__47436),
            .I(N__47127));
    ClkMux I__11135 (
            .O(N__47435),
            .I(N__47127));
    ClkMux I__11134 (
            .O(N__47434),
            .I(N__47127));
    ClkMux I__11133 (
            .O(N__47433),
            .I(N__47127));
    ClkMux I__11132 (
            .O(N__47432),
            .I(N__47127));
    ClkMux I__11131 (
            .O(N__47431),
            .I(N__47127));
    ClkMux I__11130 (
            .O(N__47430),
            .I(N__47127));
    ClkMux I__11129 (
            .O(N__47429),
            .I(N__47127));
    ClkMux I__11128 (
            .O(N__47428),
            .I(N__47127));
    ClkMux I__11127 (
            .O(N__47427),
            .I(N__47127));
    ClkMux I__11126 (
            .O(N__47426),
            .I(N__47127));
    ClkMux I__11125 (
            .O(N__47425),
            .I(N__47127));
    ClkMux I__11124 (
            .O(N__47424),
            .I(N__47127));
    ClkMux I__11123 (
            .O(N__47423),
            .I(N__47127));
    ClkMux I__11122 (
            .O(N__47422),
            .I(N__47127));
    ClkMux I__11121 (
            .O(N__47421),
            .I(N__47127));
    ClkMux I__11120 (
            .O(N__47420),
            .I(N__47127));
    ClkMux I__11119 (
            .O(N__47419),
            .I(N__47127));
    ClkMux I__11118 (
            .O(N__47418),
            .I(N__47127));
    ClkMux I__11117 (
            .O(N__47417),
            .I(N__47127));
    ClkMux I__11116 (
            .O(N__47416),
            .I(N__47127));
    Glb2LocalMux I__11115 (
            .O(N__47413),
            .I(N__47127));
    ClkMux I__11114 (
            .O(N__47412),
            .I(N__47127));
    GlobalMux I__11113 (
            .O(N__47127),
            .I(clock_output_0));
    InMux I__11112 (
            .O(N__47124),
            .I(N__47118));
    InMux I__11111 (
            .O(N__47123),
            .I(N__47115));
    InMux I__11110 (
            .O(N__47122),
            .I(N__47112));
    InMux I__11109 (
            .O(N__47121),
            .I(N__47109));
    LocalMux I__11108 (
            .O(N__47118),
            .I(N__47106));
    LocalMux I__11107 (
            .O(N__47115),
            .I(N__47103));
    LocalMux I__11106 (
            .O(N__47112),
            .I(N__47100));
    LocalMux I__11105 (
            .O(N__47109),
            .I(N__47095));
    Glb2LocalMux I__11104 (
            .O(N__47106),
            .I(N__46662));
    Glb2LocalMux I__11103 (
            .O(N__47103),
            .I(N__46662));
    Glb2LocalMux I__11102 (
            .O(N__47100),
            .I(N__46662));
    SRMux I__11101 (
            .O(N__47099),
            .I(N__46662));
    SRMux I__11100 (
            .O(N__47098),
            .I(N__46662));
    Glb2LocalMux I__11099 (
            .O(N__47095),
            .I(N__46662));
    SRMux I__11098 (
            .O(N__47094),
            .I(N__46662));
    SRMux I__11097 (
            .O(N__47093),
            .I(N__46662));
    SRMux I__11096 (
            .O(N__47092),
            .I(N__46662));
    SRMux I__11095 (
            .O(N__47091),
            .I(N__46662));
    SRMux I__11094 (
            .O(N__47090),
            .I(N__46662));
    SRMux I__11093 (
            .O(N__47089),
            .I(N__46662));
    SRMux I__11092 (
            .O(N__47088),
            .I(N__46662));
    SRMux I__11091 (
            .O(N__47087),
            .I(N__46662));
    SRMux I__11090 (
            .O(N__47086),
            .I(N__46662));
    SRMux I__11089 (
            .O(N__47085),
            .I(N__46662));
    SRMux I__11088 (
            .O(N__47084),
            .I(N__46662));
    SRMux I__11087 (
            .O(N__47083),
            .I(N__46662));
    SRMux I__11086 (
            .O(N__47082),
            .I(N__46662));
    SRMux I__11085 (
            .O(N__47081),
            .I(N__46662));
    SRMux I__11084 (
            .O(N__47080),
            .I(N__46662));
    SRMux I__11083 (
            .O(N__47079),
            .I(N__46662));
    SRMux I__11082 (
            .O(N__47078),
            .I(N__46662));
    SRMux I__11081 (
            .O(N__47077),
            .I(N__46662));
    SRMux I__11080 (
            .O(N__47076),
            .I(N__46662));
    SRMux I__11079 (
            .O(N__47075),
            .I(N__46662));
    SRMux I__11078 (
            .O(N__47074),
            .I(N__46662));
    SRMux I__11077 (
            .O(N__47073),
            .I(N__46662));
    SRMux I__11076 (
            .O(N__47072),
            .I(N__46662));
    SRMux I__11075 (
            .O(N__47071),
            .I(N__46662));
    SRMux I__11074 (
            .O(N__47070),
            .I(N__46662));
    SRMux I__11073 (
            .O(N__47069),
            .I(N__46662));
    SRMux I__11072 (
            .O(N__47068),
            .I(N__46662));
    SRMux I__11071 (
            .O(N__47067),
            .I(N__46662));
    SRMux I__11070 (
            .O(N__47066),
            .I(N__46662));
    SRMux I__11069 (
            .O(N__47065),
            .I(N__46662));
    SRMux I__11068 (
            .O(N__47064),
            .I(N__46662));
    SRMux I__11067 (
            .O(N__47063),
            .I(N__46662));
    SRMux I__11066 (
            .O(N__47062),
            .I(N__46662));
    SRMux I__11065 (
            .O(N__47061),
            .I(N__46662));
    SRMux I__11064 (
            .O(N__47060),
            .I(N__46662));
    SRMux I__11063 (
            .O(N__47059),
            .I(N__46662));
    SRMux I__11062 (
            .O(N__47058),
            .I(N__46662));
    SRMux I__11061 (
            .O(N__47057),
            .I(N__46662));
    SRMux I__11060 (
            .O(N__47056),
            .I(N__46662));
    SRMux I__11059 (
            .O(N__47055),
            .I(N__46662));
    SRMux I__11058 (
            .O(N__47054),
            .I(N__46662));
    SRMux I__11057 (
            .O(N__47053),
            .I(N__46662));
    SRMux I__11056 (
            .O(N__47052),
            .I(N__46662));
    SRMux I__11055 (
            .O(N__47051),
            .I(N__46662));
    SRMux I__11054 (
            .O(N__47050),
            .I(N__46662));
    SRMux I__11053 (
            .O(N__47049),
            .I(N__46662));
    SRMux I__11052 (
            .O(N__47048),
            .I(N__46662));
    SRMux I__11051 (
            .O(N__47047),
            .I(N__46662));
    SRMux I__11050 (
            .O(N__47046),
            .I(N__46662));
    SRMux I__11049 (
            .O(N__47045),
            .I(N__46662));
    SRMux I__11048 (
            .O(N__47044),
            .I(N__46662));
    SRMux I__11047 (
            .O(N__47043),
            .I(N__46662));
    SRMux I__11046 (
            .O(N__47042),
            .I(N__46662));
    SRMux I__11045 (
            .O(N__47041),
            .I(N__46662));
    SRMux I__11044 (
            .O(N__47040),
            .I(N__46662));
    SRMux I__11043 (
            .O(N__47039),
            .I(N__46662));
    SRMux I__11042 (
            .O(N__47038),
            .I(N__46662));
    SRMux I__11041 (
            .O(N__47037),
            .I(N__46662));
    SRMux I__11040 (
            .O(N__47036),
            .I(N__46662));
    SRMux I__11039 (
            .O(N__47035),
            .I(N__46662));
    SRMux I__11038 (
            .O(N__47034),
            .I(N__46662));
    SRMux I__11037 (
            .O(N__47033),
            .I(N__46662));
    SRMux I__11036 (
            .O(N__47032),
            .I(N__46662));
    SRMux I__11035 (
            .O(N__47031),
            .I(N__46662));
    SRMux I__11034 (
            .O(N__47030),
            .I(N__46662));
    SRMux I__11033 (
            .O(N__47029),
            .I(N__46662));
    SRMux I__11032 (
            .O(N__47028),
            .I(N__46662));
    SRMux I__11031 (
            .O(N__47027),
            .I(N__46662));
    SRMux I__11030 (
            .O(N__47026),
            .I(N__46662));
    SRMux I__11029 (
            .O(N__47025),
            .I(N__46662));
    SRMux I__11028 (
            .O(N__47024),
            .I(N__46662));
    SRMux I__11027 (
            .O(N__47023),
            .I(N__46662));
    SRMux I__11026 (
            .O(N__47022),
            .I(N__46662));
    SRMux I__11025 (
            .O(N__47021),
            .I(N__46662));
    SRMux I__11024 (
            .O(N__47020),
            .I(N__46662));
    SRMux I__11023 (
            .O(N__47019),
            .I(N__46662));
    SRMux I__11022 (
            .O(N__47018),
            .I(N__46662));
    SRMux I__11021 (
            .O(N__47017),
            .I(N__46662));
    SRMux I__11020 (
            .O(N__47016),
            .I(N__46662));
    SRMux I__11019 (
            .O(N__47015),
            .I(N__46662));
    SRMux I__11018 (
            .O(N__47014),
            .I(N__46662));
    SRMux I__11017 (
            .O(N__47013),
            .I(N__46662));
    SRMux I__11016 (
            .O(N__47012),
            .I(N__46662));
    SRMux I__11015 (
            .O(N__47011),
            .I(N__46662));
    SRMux I__11014 (
            .O(N__47010),
            .I(N__46662));
    SRMux I__11013 (
            .O(N__47009),
            .I(N__46662));
    SRMux I__11012 (
            .O(N__47008),
            .I(N__46662));
    SRMux I__11011 (
            .O(N__47007),
            .I(N__46662));
    SRMux I__11010 (
            .O(N__47006),
            .I(N__46662));
    SRMux I__11009 (
            .O(N__47005),
            .I(N__46662));
    SRMux I__11008 (
            .O(N__47004),
            .I(N__46662));
    SRMux I__11007 (
            .O(N__47003),
            .I(N__46662));
    SRMux I__11006 (
            .O(N__47002),
            .I(N__46662));
    SRMux I__11005 (
            .O(N__47001),
            .I(N__46662));
    SRMux I__11004 (
            .O(N__47000),
            .I(N__46662));
    SRMux I__11003 (
            .O(N__46999),
            .I(N__46662));
    SRMux I__11002 (
            .O(N__46998),
            .I(N__46662));
    SRMux I__11001 (
            .O(N__46997),
            .I(N__46662));
    SRMux I__11000 (
            .O(N__46996),
            .I(N__46662));
    SRMux I__10999 (
            .O(N__46995),
            .I(N__46662));
    SRMux I__10998 (
            .O(N__46994),
            .I(N__46662));
    SRMux I__10997 (
            .O(N__46993),
            .I(N__46662));
    SRMux I__10996 (
            .O(N__46992),
            .I(N__46662));
    SRMux I__10995 (
            .O(N__46991),
            .I(N__46662));
    SRMux I__10994 (
            .O(N__46990),
            .I(N__46662));
    SRMux I__10993 (
            .O(N__46989),
            .I(N__46662));
    SRMux I__10992 (
            .O(N__46988),
            .I(N__46662));
    SRMux I__10991 (
            .O(N__46987),
            .I(N__46662));
    SRMux I__10990 (
            .O(N__46986),
            .I(N__46662));
    SRMux I__10989 (
            .O(N__46985),
            .I(N__46662));
    SRMux I__10988 (
            .O(N__46984),
            .I(N__46662));
    SRMux I__10987 (
            .O(N__46983),
            .I(N__46662));
    SRMux I__10986 (
            .O(N__46982),
            .I(N__46662));
    SRMux I__10985 (
            .O(N__46981),
            .I(N__46662));
    SRMux I__10984 (
            .O(N__46980),
            .I(N__46662));
    SRMux I__10983 (
            .O(N__46979),
            .I(N__46662));
    SRMux I__10982 (
            .O(N__46978),
            .I(N__46662));
    SRMux I__10981 (
            .O(N__46977),
            .I(N__46662));
    SRMux I__10980 (
            .O(N__46976),
            .I(N__46662));
    SRMux I__10979 (
            .O(N__46975),
            .I(N__46662));
    SRMux I__10978 (
            .O(N__46974),
            .I(N__46662));
    SRMux I__10977 (
            .O(N__46973),
            .I(N__46662));
    SRMux I__10976 (
            .O(N__46972),
            .I(N__46662));
    SRMux I__10975 (
            .O(N__46971),
            .I(N__46662));
    SRMux I__10974 (
            .O(N__46970),
            .I(N__46662));
    SRMux I__10973 (
            .O(N__46969),
            .I(N__46662));
    SRMux I__10972 (
            .O(N__46968),
            .I(N__46662));
    SRMux I__10971 (
            .O(N__46967),
            .I(N__46662));
    SRMux I__10970 (
            .O(N__46966),
            .I(N__46662));
    SRMux I__10969 (
            .O(N__46965),
            .I(N__46662));
    SRMux I__10968 (
            .O(N__46964),
            .I(N__46662));
    SRMux I__10967 (
            .O(N__46963),
            .I(N__46662));
    SRMux I__10966 (
            .O(N__46962),
            .I(N__46662));
    SRMux I__10965 (
            .O(N__46961),
            .I(N__46662));
    SRMux I__10964 (
            .O(N__46960),
            .I(N__46662));
    SRMux I__10963 (
            .O(N__46959),
            .I(N__46662));
    SRMux I__10962 (
            .O(N__46958),
            .I(N__46662));
    SRMux I__10961 (
            .O(N__46957),
            .I(N__46662));
    SRMux I__10960 (
            .O(N__46956),
            .I(N__46662));
    SRMux I__10959 (
            .O(N__46955),
            .I(N__46662));
    GlobalMux I__10958 (
            .O(N__46662),
            .I(N__46659));
    gio2CtrlBuf I__10957 (
            .O(N__46659),
            .I(red_c_g));
    CascadeMux I__10956 (
            .O(N__46656),
            .I(N__46652));
    InMux I__10955 (
            .O(N__46655),
            .I(N__46647));
    InMux I__10954 (
            .O(N__46652),
            .I(N__46644));
    InMux I__10953 (
            .O(N__46651),
            .I(N__46641));
    InMux I__10952 (
            .O(N__46650),
            .I(N__46638));
    LocalMux I__10951 (
            .O(N__46647),
            .I(N__46634));
    LocalMux I__10950 (
            .O(N__46644),
            .I(N__46631));
    LocalMux I__10949 (
            .O(N__46641),
            .I(N__46626));
    LocalMux I__10948 (
            .O(N__46638),
            .I(N__46626));
    InMux I__10947 (
            .O(N__46637),
            .I(N__46623));
    Span4Mux_h I__10946 (
            .O(N__46634),
            .I(N__46620));
    Span4Mux_h I__10945 (
            .O(N__46631),
            .I(N__46613));
    Span4Mux_v I__10944 (
            .O(N__46626),
            .I(N__46613));
    LocalMux I__10943 (
            .O(N__46623),
            .I(N__46613));
    Odrv4 I__10942 (
            .O(N__46620),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__10941 (
            .O(N__46613),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    CascadeMux I__10940 (
            .O(N__46608),
            .I(N__46605));
    InMux I__10939 (
            .O(N__46605),
            .I(N__46601));
    InMux I__10938 (
            .O(N__46604),
            .I(N__46598));
    LocalMux I__10937 (
            .O(N__46601),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    LocalMux I__10936 (
            .O(N__46598),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    InMux I__10935 (
            .O(N__46593),
            .I(N__46589));
    CascadeMux I__10934 (
            .O(N__46592),
            .I(N__46584));
    LocalMux I__10933 (
            .O(N__46589),
            .I(N__46581));
    InMux I__10932 (
            .O(N__46588),
            .I(N__46578));
    InMux I__10931 (
            .O(N__46587),
            .I(N__46573));
    InMux I__10930 (
            .O(N__46584),
            .I(N__46573));
    Span4Mux_v I__10929 (
            .O(N__46581),
            .I(N__46568));
    LocalMux I__10928 (
            .O(N__46578),
            .I(N__46568));
    LocalMux I__10927 (
            .O(N__46573),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__10926 (
            .O(N__46568),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__10925 (
            .O(N__46563),
            .I(N__46560));
    LocalMux I__10924 (
            .O(N__46560),
            .I(N__46555));
    InMux I__10923 (
            .O(N__46559),
            .I(N__46550));
    InMux I__10922 (
            .O(N__46558),
            .I(N__46550));
    Span4Mux_v I__10921 (
            .O(N__46555),
            .I(N__46547));
    LocalMux I__10920 (
            .O(N__46550),
            .I(N__46543));
    Sp12to4 I__10919 (
            .O(N__46547),
            .I(N__46540));
    InMux I__10918 (
            .O(N__46546),
            .I(N__46537));
    Span4Mux_v I__10917 (
            .O(N__46543),
            .I(N__46533));
    Span12Mux_h I__10916 (
            .O(N__46540),
            .I(N__46530));
    LocalMux I__10915 (
            .O(N__46537),
            .I(N__46527));
    InMux I__10914 (
            .O(N__46536),
            .I(N__46524));
    Span4Mux_h I__10913 (
            .O(N__46533),
            .I(N__46521));
    Odrv12 I__10912 (
            .O(N__46530),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv12 I__10911 (
            .O(N__46527),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__10910 (
            .O(N__46524),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv4 I__10909 (
            .O(N__46521),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    CascadeMux I__10908 (
            .O(N__46512),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24_cascade_));
    InMux I__10907 (
            .O(N__46509),
            .I(N__46506));
    LocalMux I__10906 (
            .O(N__46506),
            .I(N__46503));
    Span4Mux_v I__10905 (
            .O(N__46503),
            .I(N__46498));
    InMux I__10904 (
            .O(N__46502),
            .I(N__46493));
    InMux I__10903 (
            .O(N__46501),
            .I(N__46493));
    Sp12to4 I__10902 (
            .O(N__46498),
            .I(N__46488));
    LocalMux I__10901 (
            .O(N__46493),
            .I(N__46488));
    Span12Mux_h I__10900 (
            .O(N__46488),
            .I(N__46484));
    InMux I__10899 (
            .O(N__46487),
            .I(N__46481));
    Odrv12 I__10898 (
            .O(N__46484),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__10897 (
            .O(N__46481),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__10896 (
            .O(N__46476),
            .I(N__46470));
    InMux I__10895 (
            .O(N__46475),
            .I(N__46470));
    LocalMux I__10894 (
            .O(N__46470),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    InMux I__10893 (
            .O(N__46467),
            .I(N__46463));
    InMux I__10892 (
            .O(N__46466),
            .I(N__46460));
    LocalMux I__10891 (
            .O(N__46463),
            .I(N__46457));
    LocalMux I__10890 (
            .O(N__46460),
            .I(N__46452));
    Span4Mux_h I__10889 (
            .O(N__46457),
            .I(N__46449));
    InMux I__10888 (
            .O(N__46456),
            .I(N__46446));
    InMux I__10887 (
            .O(N__46455),
            .I(N__46443));
    Span4Mux_v I__10886 (
            .O(N__46452),
            .I(N__46440));
    Sp12to4 I__10885 (
            .O(N__46449),
            .I(N__46435));
    LocalMux I__10884 (
            .O(N__46446),
            .I(N__46435));
    LocalMux I__10883 (
            .O(N__46443),
            .I(N__46430));
    Sp12to4 I__10882 (
            .O(N__46440),
            .I(N__46425));
    Span12Mux_s8_v I__10881 (
            .O(N__46435),
            .I(N__46425));
    InMux I__10880 (
            .O(N__46434),
            .I(N__46420));
    InMux I__10879 (
            .O(N__46433),
            .I(N__46420));
    Odrv12 I__10878 (
            .O(N__46430),
            .I(phase_controller_inst1_state_4));
    Odrv12 I__10877 (
            .O(N__46425),
            .I(phase_controller_inst1_state_4));
    LocalMux I__10876 (
            .O(N__46420),
            .I(phase_controller_inst1_state_4));
    InMux I__10875 (
            .O(N__46413),
            .I(N__46410));
    LocalMux I__10874 (
            .O(N__46410),
            .I(N__46407));
    Span4Mux_v I__10873 (
            .O(N__46407),
            .I(N__46404));
    Span4Mux_h I__10872 (
            .O(N__46404),
            .I(N__46401));
    Odrv4 I__10871 (
            .O(N__46401),
            .I(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ));
    InMux I__10870 (
            .O(N__46398),
            .I(N__46395));
    LocalMux I__10869 (
            .O(N__46395),
            .I(N__46392));
    Span4Mux_h I__10868 (
            .O(N__46392),
            .I(N__46389));
    Span4Mux_h I__10867 (
            .O(N__46389),
            .I(N__46385));
    InMux I__10866 (
            .O(N__46388),
            .I(N__46382));
    Odrv4 I__10865 (
            .O(N__46385),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    LocalMux I__10864 (
            .O(N__46382),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    CascadeMux I__10863 (
            .O(N__46377),
            .I(N__46374));
    InMux I__10862 (
            .O(N__46374),
            .I(N__46369));
    InMux I__10861 (
            .O(N__46373),
            .I(N__46366));
    InMux I__10860 (
            .O(N__46372),
            .I(N__46363));
    LocalMux I__10859 (
            .O(N__46369),
            .I(N__46360));
    LocalMux I__10858 (
            .O(N__46366),
            .I(N__46357));
    LocalMux I__10857 (
            .O(N__46363),
            .I(N__46354));
    Span4Mux_h I__10856 (
            .O(N__46360),
            .I(N__46350));
    Span4Mux_h I__10855 (
            .O(N__46357),
            .I(N__46345));
    Span4Mux_v I__10854 (
            .O(N__46354),
            .I(N__46345));
    InMux I__10853 (
            .O(N__46353),
            .I(N__46342));
    Odrv4 I__10852 (
            .O(N__46350),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__10851 (
            .O(N__46345),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__10850 (
            .O(N__46342),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__10849 (
            .O(N__46335),
            .I(N__46332));
    LocalMux I__10848 (
            .O(N__46332),
            .I(N__46329));
    Span4Mux_h I__10847 (
            .O(N__46329),
            .I(N__46326));
    Odrv4 I__10846 (
            .O(N__46326),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    CascadeMux I__10845 (
            .O(N__46323),
            .I(N__46320));
    InMux I__10844 (
            .O(N__46320),
            .I(N__46315));
    InMux I__10843 (
            .O(N__46319),
            .I(N__46312));
    InMux I__10842 (
            .O(N__46318),
            .I(N__46309));
    LocalMux I__10841 (
            .O(N__46315),
            .I(N__46304));
    LocalMux I__10840 (
            .O(N__46312),
            .I(N__46304));
    LocalMux I__10839 (
            .O(N__46309),
            .I(N__46301));
    Span4Mux_v I__10838 (
            .O(N__46304),
            .I(N__46295));
    Span4Mux_v I__10837 (
            .O(N__46301),
            .I(N__46295));
    InMux I__10836 (
            .O(N__46300),
            .I(N__46292));
    Odrv4 I__10835 (
            .O(N__46295),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__10834 (
            .O(N__46292),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__10833 (
            .O(N__46287),
            .I(N__46284));
    LocalMux I__10832 (
            .O(N__46284),
            .I(N__46281));
    Span4Mux_h I__10831 (
            .O(N__46281),
            .I(N__46278));
    Odrv4 I__10830 (
            .O(N__46278),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    CascadeMux I__10829 (
            .O(N__46275),
            .I(N__46272));
    InMux I__10828 (
            .O(N__46272),
            .I(N__46268));
    InMux I__10827 (
            .O(N__46271),
            .I(N__46264));
    LocalMux I__10826 (
            .O(N__46268),
            .I(N__46261));
    InMux I__10825 (
            .O(N__46267),
            .I(N__46258));
    LocalMux I__10824 (
            .O(N__46264),
            .I(N__46255));
    Span4Mux_v I__10823 (
            .O(N__46261),
            .I(N__46252));
    LocalMux I__10822 (
            .O(N__46258),
            .I(N__46249));
    Span4Mux_h I__10821 (
            .O(N__46255),
            .I(N__46245));
    Span4Mux_h I__10820 (
            .O(N__46252),
            .I(N__46240));
    Span4Mux_v I__10819 (
            .O(N__46249),
            .I(N__46240));
    InMux I__10818 (
            .O(N__46248),
            .I(N__46237));
    Odrv4 I__10817 (
            .O(N__46245),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__10816 (
            .O(N__46240),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__10815 (
            .O(N__46237),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__10814 (
            .O(N__46230),
            .I(N__46227));
    LocalMux I__10813 (
            .O(N__46227),
            .I(N__46224));
    Span4Mux_h I__10812 (
            .O(N__46224),
            .I(N__46221));
    Odrv4 I__10811 (
            .O(N__46221),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__10810 (
            .O(N__46218),
            .I(N__46214));
    InMux I__10809 (
            .O(N__46217),
            .I(N__46211));
    LocalMux I__10808 (
            .O(N__46214),
            .I(N__46205));
    LocalMux I__10807 (
            .O(N__46211),
            .I(N__46205));
    InMux I__10806 (
            .O(N__46210),
            .I(N__46201));
    Span4Mux_v I__10805 (
            .O(N__46205),
            .I(N__46198));
    InMux I__10804 (
            .O(N__46204),
            .I(N__46195));
    LocalMux I__10803 (
            .O(N__46201),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__10802 (
            .O(N__46198),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__10801 (
            .O(N__46195),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__10800 (
            .O(N__46188),
            .I(N__46185));
    LocalMux I__10799 (
            .O(N__46185),
            .I(N__46182));
    Span4Mux_h I__10798 (
            .O(N__46182),
            .I(N__46179));
    Odrv4 I__10797 (
            .O(N__46179),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__10796 (
            .O(N__46176),
            .I(N__46173));
    LocalMux I__10795 (
            .O(N__46173),
            .I(N__46168));
    InMux I__10794 (
            .O(N__46172),
            .I(N__46165));
    InMux I__10793 (
            .O(N__46171),
            .I(N__46162));
    Span12Mux_s11_v I__10792 (
            .O(N__46168),
            .I(N__46157));
    LocalMux I__10791 (
            .O(N__46165),
            .I(N__46157));
    LocalMux I__10790 (
            .O(N__46162),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    Odrv12 I__10789 (
            .O(N__46157),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    InMux I__10788 (
            .O(N__46152),
            .I(N__46149));
    LocalMux I__10787 (
            .O(N__46149),
            .I(N__46143));
    InMux I__10786 (
            .O(N__46148),
            .I(N__46140));
    CascadeMux I__10785 (
            .O(N__46147),
            .I(N__46137));
    InMux I__10784 (
            .O(N__46146),
            .I(N__46134));
    Span4Mux_h I__10783 (
            .O(N__46143),
            .I(N__46131));
    LocalMux I__10782 (
            .O(N__46140),
            .I(N__46128));
    InMux I__10781 (
            .O(N__46137),
            .I(N__46125));
    LocalMux I__10780 (
            .O(N__46134),
            .I(N__46122));
    Span4Mux_h I__10779 (
            .O(N__46131),
            .I(N__46117));
    Span4Mux_v I__10778 (
            .O(N__46128),
            .I(N__46117));
    LocalMux I__10777 (
            .O(N__46125),
            .I(N__46114));
    Odrv12 I__10776 (
            .O(N__46122),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv4 I__10775 (
            .O(N__46117),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv4 I__10774 (
            .O(N__46114),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__10773 (
            .O(N__46107),
            .I(N__46104));
    LocalMux I__10772 (
            .O(N__46104),
            .I(N__46101));
    Span4Mux_h I__10771 (
            .O(N__46101),
            .I(N__46098));
    Odrv4 I__10770 (
            .O(N__46098),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    InMux I__10769 (
            .O(N__46095),
            .I(N__46092));
    LocalMux I__10768 (
            .O(N__46092),
            .I(N__46089));
    Span4Mux_h I__10767 (
            .O(N__46089),
            .I(N__46086));
    Odrv4 I__10766 (
            .O(N__46086),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CEMux I__10765 (
            .O(N__46083),
            .I(N__46059));
    CEMux I__10764 (
            .O(N__46082),
            .I(N__46059));
    CEMux I__10763 (
            .O(N__46081),
            .I(N__46059));
    CEMux I__10762 (
            .O(N__46080),
            .I(N__46059));
    CEMux I__10761 (
            .O(N__46079),
            .I(N__46059));
    CEMux I__10760 (
            .O(N__46078),
            .I(N__46059));
    CEMux I__10759 (
            .O(N__46077),
            .I(N__46059));
    CEMux I__10758 (
            .O(N__46076),
            .I(N__46059));
    GlobalMux I__10757 (
            .O(N__46059),
            .I(N__46056));
    gio2CtrlBuf I__10756 (
            .O(N__46056),
            .I(\phase_controller_inst2.stoper_tr.un1_start_g ));
    InMux I__10755 (
            .O(N__46053),
            .I(N__46050));
    LocalMux I__10754 (
            .O(N__46050),
            .I(N__46047));
    Odrv12 I__10753 (
            .O(N__46047),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ));
    InMux I__10752 (
            .O(N__46044),
            .I(N__46038));
    InMux I__10751 (
            .O(N__46043),
            .I(N__46038));
    LocalMux I__10750 (
            .O(N__46038),
            .I(N__46034));
    InMux I__10749 (
            .O(N__46037),
            .I(N__46031));
    Span4Mux_h I__10748 (
            .O(N__46034),
            .I(N__46028));
    LocalMux I__10747 (
            .O(N__46031),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__10746 (
            .O(N__46028),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    CascadeMux I__10745 (
            .O(N__46023),
            .I(N__46019));
    InMux I__10744 (
            .O(N__46022),
            .I(N__46014));
    InMux I__10743 (
            .O(N__46019),
            .I(N__46014));
    LocalMux I__10742 (
            .O(N__46014),
            .I(N__46010));
    InMux I__10741 (
            .O(N__46013),
            .I(N__46007));
    Span4Mux_h I__10740 (
            .O(N__46010),
            .I(N__46004));
    LocalMux I__10739 (
            .O(N__46007),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__10738 (
            .O(N__46004),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__10737 (
            .O(N__45999),
            .I(N__45993));
    InMux I__10736 (
            .O(N__45998),
            .I(N__45993));
    LocalMux I__10735 (
            .O(N__45993),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ));
    CascadeMux I__10734 (
            .O(N__45990),
            .I(N__45987));
    InMux I__10733 (
            .O(N__45987),
            .I(N__45984));
    LocalMux I__10732 (
            .O(N__45984),
            .I(N__45981));
    Odrv12 I__10731 (
            .O(N__45981),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt28 ));
    CascadeMux I__10730 (
            .O(N__45978),
            .I(N__45974));
    InMux I__10729 (
            .O(N__45977),
            .I(N__45971));
    InMux I__10728 (
            .O(N__45974),
            .I(N__45968));
    LocalMux I__10727 (
            .O(N__45971),
            .I(N__45963));
    LocalMux I__10726 (
            .O(N__45968),
            .I(N__45963));
    Span4Mux_v I__10725 (
            .O(N__45963),
            .I(N__45960));
    Odrv4 I__10724 (
            .O(N__45960),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    InMux I__10723 (
            .O(N__45957),
            .I(N__45954));
    LocalMux I__10722 (
            .O(N__45954),
            .I(N__45950));
    InMux I__10721 (
            .O(N__45953),
            .I(N__45946));
    Span4Mux_h I__10720 (
            .O(N__45950),
            .I(N__45943));
    InMux I__10719 (
            .O(N__45949),
            .I(N__45940));
    LocalMux I__10718 (
            .O(N__45946),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__10717 (
            .O(N__45943),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__10716 (
            .O(N__45940),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    CascadeMux I__10715 (
            .O(N__45933),
            .I(N__45930));
    InMux I__10714 (
            .O(N__45930),
            .I(N__45927));
    LocalMux I__10713 (
            .O(N__45927),
            .I(N__45922));
    InMux I__10712 (
            .O(N__45926),
            .I(N__45919));
    InMux I__10711 (
            .O(N__45925),
            .I(N__45916));
    Span4Mux_v I__10710 (
            .O(N__45922),
            .I(N__45913));
    LocalMux I__10709 (
            .O(N__45919),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__10708 (
            .O(N__45916),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv4 I__10707 (
            .O(N__45913),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__10706 (
            .O(N__45906),
            .I(N__45902));
    InMux I__10705 (
            .O(N__45905),
            .I(N__45899));
    LocalMux I__10704 (
            .O(N__45902),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    LocalMux I__10703 (
            .O(N__45899),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    CascadeMux I__10702 (
            .O(N__45894),
            .I(N__45891));
    InMux I__10701 (
            .O(N__45891),
            .I(N__45888));
    LocalMux I__10700 (
            .O(N__45888),
            .I(N__45885));
    Odrv12 I__10699 (
            .O(N__45885),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt26 ));
    CascadeMux I__10698 (
            .O(N__45882),
            .I(N__45879));
    InMux I__10697 (
            .O(N__45879),
            .I(N__45876));
    LocalMux I__10696 (
            .O(N__45876),
            .I(N__45873));
    Span4Mux_v I__10695 (
            .O(N__45873),
            .I(N__45870));
    Span4Mux_h I__10694 (
            .O(N__45870),
            .I(N__45867));
    Odrv4 I__10693 (
            .O(N__45867),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt24 ));
    CascadeMux I__10692 (
            .O(N__45864),
            .I(N__45860));
    InMux I__10691 (
            .O(N__45863),
            .I(N__45855));
    InMux I__10690 (
            .O(N__45860),
            .I(N__45855));
    LocalMux I__10689 (
            .O(N__45855),
            .I(N__45851));
    InMux I__10688 (
            .O(N__45854),
            .I(N__45848));
    Span4Mux_h I__10687 (
            .O(N__45851),
            .I(N__45845));
    LocalMux I__10686 (
            .O(N__45848),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__10685 (
            .O(N__45845),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    CascadeMux I__10684 (
            .O(N__45840),
            .I(N__45836));
    InMux I__10683 (
            .O(N__45839),
            .I(N__45832));
    InMux I__10682 (
            .O(N__45836),
            .I(N__45827));
    InMux I__10681 (
            .O(N__45835),
            .I(N__45827));
    LocalMux I__10680 (
            .O(N__45832),
            .I(N__45822));
    LocalMux I__10679 (
            .O(N__45827),
            .I(N__45822));
    Odrv4 I__10678 (
            .O(N__45822),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__10677 (
            .O(N__45819),
            .I(N__45816));
    LocalMux I__10676 (
            .O(N__45816),
            .I(N__45813));
    Span4Mux_v I__10675 (
            .O(N__45813),
            .I(N__45810));
    Span4Mux_h I__10674 (
            .O(N__45810),
            .I(N__45807));
    Odrv4 I__10673 (
            .O(N__45807),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ));
    InMux I__10672 (
            .O(N__45804),
            .I(N__45801));
    LocalMux I__10671 (
            .O(N__45801),
            .I(N__45797));
    InMux I__10670 (
            .O(N__45800),
            .I(N__45794));
    Odrv4 I__10669 (
            .O(N__45797),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    LocalMux I__10668 (
            .O(N__45794),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    CascadeMux I__10667 (
            .O(N__45789),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_));
    InMux I__10666 (
            .O(N__45786),
            .I(N__45783));
    LocalMux I__10665 (
            .O(N__45783),
            .I(N__45778));
    InMux I__10664 (
            .O(N__45782),
            .I(N__45773));
    InMux I__10663 (
            .O(N__45781),
            .I(N__45773));
    Span4Mux_h I__10662 (
            .O(N__45778),
            .I(N__45768));
    LocalMux I__10661 (
            .O(N__45773),
            .I(N__45768));
    Span4Mux_v I__10660 (
            .O(N__45768),
            .I(N__45764));
    CascadeMux I__10659 (
            .O(N__45767),
            .I(N__45761));
    Span4Mux_h I__10658 (
            .O(N__45764),
            .I(N__45758));
    InMux I__10657 (
            .O(N__45761),
            .I(N__45755));
    Odrv4 I__10656 (
            .O(N__45758),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__10655 (
            .O(N__45755),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__10654 (
            .O(N__45750),
            .I(N__45744));
    InMux I__10653 (
            .O(N__45749),
            .I(N__45744));
    LocalMux I__10652 (
            .O(N__45744),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ));
    InMux I__10651 (
            .O(N__45741),
            .I(N__45738));
    LocalMux I__10650 (
            .O(N__45738),
            .I(N__45734));
    InMux I__10649 (
            .O(N__45737),
            .I(N__45731));
    Odrv4 I__10648 (
            .O(N__45734),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    LocalMux I__10647 (
            .O(N__45731),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__10646 (
            .O(N__45726),
            .I(N__45720));
    InMux I__10645 (
            .O(N__45725),
            .I(N__45720));
    LocalMux I__10644 (
            .O(N__45720),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    InMux I__10643 (
            .O(N__45717),
            .I(N__45711));
    InMux I__10642 (
            .O(N__45716),
            .I(N__45711));
    LocalMux I__10641 (
            .O(N__45711),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    InMux I__10640 (
            .O(N__45708),
            .I(N__45702));
    InMux I__10639 (
            .O(N__45707),
            .I(N__45702));
    LocalMux I__10638 (
            .O(N__45702),
            .I(N__45699));
    Odrv4 I__10637 (
            .O(N__45699),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    CascadeMux I__10636 (
            .O(N__45696),
            .I(N__45693));
    InMux I__10635 (
            .O(N__45693),
            .I(N__45687));
    InMux I__10634 (
            .O(N__45692),
            .I(N__45687));
    LocalMux I__10633 (
            .O(N__45687),
            .I(N__45684));
    Odrv4 I__10632 (
            .O(N__45684),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    CascadeMux I__10631 (
            .O(N__45681),
            .I(N__45678));
    InMux I__10630 (
            .O(N__45678),
            .I(N__45672));
    InMux I__10629 (
            .O(N__45677),
            .I(N__45672));
    LocalMux I__10628 (
            .O(N__45672),
            .I(N__45669));
    Odrv4 I__10627 (
            .O(N__45669),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    InMux I__10626 (
            .O(N__45666),
            .I(N__45662));
    InMux I__10625 (
            .O(N__45665),
            .I(N__45659));
    LocalMux I__10624 (
            .O(N__45662),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    LocalMux I__10623 (
            .O(N__45659),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    CascadeMux I__10622 (
            .O(N__45654),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_));
    InMux I__10621 (
            .O(N__45651),
            .I(N__45645));
    InMux I__10620 (
            .O(N__45650),
            .I(N__45640));
    InMux I__10619 (
            .O(N__45649),
            .I(N__45640));
    InMux I__10618 (
            .O(N__45648),
            .I(N__45637));
    LocalMux I__10617 (
            .O(N__45645),
            .I(N__45632));
    LocalMux I__10616 (
            .O(N__45640),
            .I(N__45632));
    LocalMux I__10615 (
            .O(N__45637),
            .I(N__45629));
    Span4Mux_v I__10614 (
            .O(N__45632),
            .I(N__45626));
    Span4Mux_h I__10613 (
            .O(N__45629),
            .I(N__45623));
    Span4Mux_h I__10612 (
            .O(N__45626),
            .I(N__45620));
    Span4Mux_h I__10611 (
            .O(N__45623),
            .I(N__45617));
    Odrv4 I__10610 (
            .O(N__45620),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__10609 (
            .O(N__45617),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__10608 (
            .O(N__45612),
            .I(N__45608));
    InMux I__10607 (
            .O(N__45611),
            .I(N__45605));
    LocalMux I__10606 (
            .O(N__45608),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    LocalMux I__10605 (
            .O(N__45605),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    CascadeMux I__10604 (
            .O(N__45600),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_));
    InMux I__10603 (
            .O(N__45597),
            .I(N__45592));
    InMux I__10602 (
            .O(N__45596),
            .I(N__45587));
    InMux I__10601 (
            .O(N__45595),
            .I(N__45587));
    LocalMux I__10600 (
            .O(N__45592),
            .I(N__45581));
    LocalMux I__10599 (
            .O(N__45587),
            .I(N__45581));
    InMux I__10598 (
            .O(N__45586),
            .I(N__45578));
    Span4Mux_v I__10597 (
            .O(N__45581),
            .I(N__45575));
    LocalMux I__10596 (
            .O(N__45578),
            .I(N__45572));
    Span4Mux_h I__10595 (
            .O(N__45575),
            .I(N__45569));
    Span12Mux_h I__10594 (
            .O(N__45572),
            .I(N__45566));
    Odrv4 I__10593 (
            .O(N__45569),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv12 I__10592 (
            .O(N__45566),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__10591 (
            .O(N__45561),
            .I(N__45558));
    LocalMux I__10590 (
            .O(N__45558),
            .I(N__45554));
    InMux I__10589 (
            .O(N__45557),
            .I(N__45551));
    Odrv4 I__10588 (
            .O(N__45554),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    LocalMux I__10587 (
            .O(N__45551),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    CascadeMux I__10586 (
            .O(N__45546),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_));
    InMux I__10585 (
            .O(N__45543),
            .I(N__45538));
    InMux I__10584 (
            .O(N__45542),
            .I(N__45533));
    InMux I__10583 (
            .O(N__45541),
            .I(N__45533));
    LocalMux I__10582 (
            .O(N__45538),
            .I(N__45530));
    LocalMux I__10581 (
            .O(N__45533),
            .I(N__45527));
    Span4Mux_h I__10580 (
            .O(N__45530),
            .I(N__45524));
    Span4Mux_h I__10579 (
            .O(N__45527),
            .I(N__45521));
    Span4Mux_h I__10578 (
            .O(N__45524),
            .I(N__45517));
    Span4Mux_h I__10577 (
            .O(N__45521),
            .I(N__45514));
    InMux I__10576 (
            .O(N__45520),
            .I(N__45511));
    Odrv4 I__10575 (
            .O(N__45517),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv4 I__10574 (
            .O(N__45514),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    LocalMux I__10573 (
            .O(N__45511),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__10572 (
            .O(N__45504),
            .I(N__45501));
    LocalMux I__10571 (
            .O(N__45501),
            .I(N__45498));
    Odrv4 I__10570 (
            .O(N__45498),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ));
    InMux I__10569 (
            .O(N__45495),
            .I(N__45490));
    InMux I__10568 (
            .O(N__45494),
            .I(N__45485));
    InMux I__10567 (
            .O(N__45493),
            .I(N__45485));
    LocalMux I__10566 (
            .O(N__45490),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__10565 (
            .O(N__45485),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    CascadeMux I__10564 (
            .O(N__45480),
            .I(N__45475));
    InMux I__10563 (
            .O(N__45479),
            .I(N__45472));
    InMux I__10562 (
            .O(N__45478),
            .I(N__45467));
    InMux I__10561 (
            .O(N__45475),
            .I(N__45467));
    LocalMux I__10560 (
            .O(N__45472),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__10559 (
            .O(N__45467),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__10558 (
            .O(N__45462),
            .I(N__45456));
    InMux I__10557 (
            .O(N__45461),
            .I(N__45456));
    LocalMux I__10556 (
            .O(N__45456),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ));
    CascadeMux I__10555 (
            .O(N__45453),
            .I(N__45450));
    InMux I__10554 (
            .O(N__45450),
            .I(N__45447));
    LocalMux I__10553 (
            .O(N__45447),
            .I(N__45444));
    Odrv4 I__10552 (
            .O(N__45444),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt26 ));
    InMux I__10551 (
            .O(N__45441),
            .I(N__45438));
    LocalMux I__10550 (
            .O(N__45438),
            .I(N__45435));
    Span4Mux_v I__10549 (
            .O(N__45435),
            .I(N__45432));
    Odrv4 I__10548 (
            .O(N__45432),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt28 ));
    CascadeMux I__10547 (
            .O(N__45429),
            .I(N__45424));
    InMux I__10546 (
            .O(N__45428),
            .I(N__45421));
    InMux I__10545 (
            .O(N__45427),
            .I(N__45416));
    InMux I__10544 (
            .O(N__45424),
            .I(N__45416));
    LocalMux I__10543 (
            .O(N__45421),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__10542 (
            .O(N__45416),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    CascadeMux I__10541 (
            .O(N__45411),
            .I(N__45406));
    InMux I__10540 (
            .O(N__45410),
            .I(N__45403));
    InMux I__10539 (
            .O(N__45409),
            .I(N__45398));
    InMux I__10538 (
            .O(N__45406),
            .I(N__45398));
    LocalMux I__10537 (
            .O(N__45403),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__10536 (
            .O(N__45398),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    CascadeMux I__10535 (
            .O(N__45393),
            .I(N__45390));
    InMux I__10534 (
            .O(N__45390),
            .I(N__45387));
    LocalMux I__10533 (
            .O(N__45387),
            .I(N__45384));
    Span4Mux_v I__10532 (
            .O(N__45384),
            .I(N__45381));
    Odrv4 I__10531 (
            .O(N__45381),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ));
    InMux I__10530 (
            .O(N__45378),
            .I(N__45374));
    InMux I__10529 (
            .O(N__45377),
            .I(N__45371));
    LocalMux I__10528 (
            .O(N__45374),
            .I(N__45364));
    LocalMux I__10527 (
            .O(N__45371),
            .I(N__45364));
    InMux I__10526 (
            .O(N__45370),
            .I(N__45361));
    InMux I__10525 (
            .O(N__45369),
            .I(N__45358));
    Span12Mux_h I__10524 (
            .O(N__45364),
            .I(N__45355));
    LocalMux I__10523 (
            .O(N__45361),
            .I(N__45350));
    LocalMux I__10522 (
            .O(N__45358),
            .I(N__45350));
    Odrv12 I__10521 (
            .O(N__45355),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv12 I__10520 (
            .O(N__45350),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__10519 (
            .O(N__45345),
            .I(N__45341));
    InMux I__10518 (
            .O(N__45344),
            .I(N__45337));
    LocalMux I__10517 (
            .O(N__45341),
            .I(N__45334));
    InMux I__10516 (
            .O(N__45340),
            .I(N__45331));
    LocalMux I__10515 (
            .O(N__45337),
            .I(N__45326));
    Span4Mux_h I__10514 (
            .O(N__45334),
            .I(N__45326));
    LocalMux I__10513 (
            .O(N__45331),
            .I(N__45323));
    Odrv4 I__10512 (
            .O(N__45326),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv12 I__10511 (
            .O(N__45323),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    InMux I__10510 (
            .O(N__45318),
            .I(N__45313));
    InMux I__10509 (
            .O(N__45317),
            .I(N__45310));
    InMux I__10508 (
            .O(N__45316),
            .I(N__45307));
    LocalMux I__10507 (
            .O(N__45313),
            .I(N__45302));
    LocalMux I__10506 (
            .O(N__45310),
            .I(N__45302));
    LocalMux I__10505 (
            .O(N__45307),
            .I(N__45298));
    Span4Mux_v I__10504 (
            .O(N__45302),
            .I(N__45295));
    InMux I__10503 (
            .O(N__45301),
            .I(N__45292));
    Span4Mux_h I__10502 (
            .O(N__45298),
            .I(N__45289));
    Span4Mux_h I__10501 (
            .O(N__45295),
            .I(N__45284));
    LocalMux I__10500 (
            .O(N__45292),
            .I(N__45284));
    Odrv4 I__10499 (
            .O(N__45289),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv4 I__10498 (
            .O(N__45284),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__10497 (
            .O(N__45279),
            .I(N__45276));
    LocalMux I__10496 (
            .O(N__45276),
            .I(N__45272));
    InMux I__10495 (
            .O(N__45275),
            .I(N__45268));
    Span4Mux_h I__10494 (
            .O(N__45272),
            .I(N__45265));
    InMux I__10493 (
            .O(N__45271),
            .I(N__45262));
    LocalMux I__10492 (
            .O(N__45268),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    Odrv4 I__10491 (
            .O(N__45265),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    LocalMux I__10490 (
            .O(N__45262),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    InMux I__10489 (
            .O(N__45255),
            .I(N__45252));
    LocalMux I__10488 (
            .O(N__45252),
            .I(N__45249));
    Span4Mux_h I__10487 (
            .O(N__45249),
            .I(N__45246));
    Odrv4 I__10486 (
            .O(N__45246),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt20 ));
    InMux I__10485 (
            .O(N__45243),
            .I(N__45238));
    InMux I__10484 (
            .O(N__45242),
            .I(N__45233));
    InMux I__10483 (
            .O(N__45241),
            .I(N__45233));
    LocalMux I__10482 (
            .O(N__45238),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    LocalMux I__10481 (
            .O(N__45233),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    CascadeMux I__10480 (
            .O(N__45228),
            .I(N__45224));
    InMux I__10479 (
            .O(N__45227),
            .I(N__45220));
    InMux I__10478 (
            .O(N__45224),
            .I(N__45215));
    InMux I__10477 (
            .O(N__45223),
            .I(N__45215));
    LocalMux I__10476 (
            .O(N__45220),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    LocalMux I__10475 (
            .O(N__45215),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    CascadeMux I__10474 (
            .O(N__45210),
            .I(N__45207));
    InMux I__10473 (
            .O(N__45207),
            .I(N__45204));
    LocalMux I__10472 (
            .O(N__45204),
            .I(N__45201));
    Span4Mux_h I__10471 (
            .O(N__45201),
            .I(N__45198));
    Odrv4 I__10470 (
            .O(N__45198),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ));
    InMux I__10469 (
            .O(N__45195),
            .I(N__45188));
    InMux I__10468 (
            .O(N__45194),
            .I(N__45188));
    InMux I__10467 (
            .O(N__45193),
            .I(N__45185));
    LocalMux I__10466 (
            .O(N__45188),
            .I(N__45182));
    LocalMux I__10465 (
            .O(N__45185),
            .I(N__45178));
    Span4Mux_h I__10464 (
            .O(N__45182),
            .I(N__45175));
    InMux I__10463 (
            .O(N__45181),
            .I(N__45172));
    Odrv12 I__10462 (
            .O(N__45178),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv4 I__10461 (
            .O(N__45175),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__10460 (
            .O(N__45172),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__10459 (
            .O(N__45165),
            .I(N__45162));
    LocalMux I__10458 (
            .O(N__45162),
            .I(N__45159));
    Span4Mux_v I__10457 (
            .O(N__45159),
            .I(N__45155));
    InMux I__10456 (
            .O(N__45158),
            .I(N__45152));
    Odrv4 I__10455 (
            .O(N__45155),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    LocalMux I__10454 (
            .O(N__45152),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    InMux I__10453 (
            .O(N__45147),
            .I(N__45141));
    InMux I__10452 (
            .O(N__45146),
            .I(N__45141));
    LocalMux I__10451 (
            .O(N__45141),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    InMux I__10450 (
            .O(N__45138),
            .I(N__45135));
    LocalMux I__10449 (
            .O(N__45135),
            .I(N__45129));
    InMux I__10448 (
            .O(N__45134),
            .I(N__45122));
    InMux I__10447 (
            .O(N__45133),
            .I(N__45122));
    InMux I__10446 (
            .O(N__45132),
            .I(N__45122));
    Odrv12 I__10445 (
            .O(N__45129),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__10444 (
            .O(N__45122),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__10443 (
            .O(N__45117),
            .I(N__45113));
    CascadeMux I__10442 (
            .O(N__45116),
            .I(N__45110));
    LocalMux I__10441 (
            .O(N__45113),
            .I(N__45107));
    InMux I__10440 (
            .O(N__45110),
            .I(N__45104));
    Span4Mux_h I__10439 (
            .O(N__45107),
            .I(N__45101));
    LocalMux I__10438 (
            .O(N__45104),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    Odrv4 I__10437 (
            .O(N__45101),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    CascadeMux I__10436 (
            .O(N__45096),
            .I(N__45093));
    InMux I__10435 (
            .O(N__45093),
            .I(N__45087));
    InMux I__10434 (
            .O(N__45092),
            .I(N__45087));
    LocalMux I__10433 (
            .O(N__45087),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    InMux I__10432 (
            .O(N__45084),
            .I(N__45081));
    LocalMux I__10431 (
            .O(N__45081),
            .I(N__45076));
    InMux I__10430 (
            .O(N__45080),
            .I(N__45073));
    InMux I__10429 (
            .O(N__45079),
            .I(N__45070));
    Span4Mux_h I__10428 (
            .O(N__45076),
            .I(N__45065));
    LocalMux I__10427 (
            .O(N__45073),
            .I(N__45065));
    LocalMux I__10426 (
            .O(N__45070),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    Odrv4 I__10425 (
            .O(N__45065),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    InMux I__10424 (
            .O(N__45060),
            .I(N__45057));
    LocalMux I__10423 (
            .O(N__45057),
            .I(N__45053));
    InMux I__10422 (
            .O(N__45056),
            .I(N__45048));
    Span4Mux_v I__10421 (
            .O(N__45053),
            .I(N__45045));
    InMux I__10420 (
            .O(N__45052),
            .I(N__45040));
    InMux I__10419 (
            .O(N__45051),
            .I(N__45040));
    LocalMux I__10418 (
            .O(N__45048),
            .I(N__45037));
    Sp12to4 I__10417 (
            .O(N__45045),
            .I(N__45032));
    LocalMux I__10416 (
            .O(N__45040),
            .I(N__45032));
    Odrv4 I__10415 (
            .O(N__45037),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv12 I__10414 (
            .O(N__45032),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    CascadeMux I__10413 (
            .O(N__45027),
            .I(N__45024));
    InMux I__10412 (
            .O(N__45024),
            .I(N__45021));
    LocalMux I__10411 (
            .O(N__45021),
            .I(N__45018));
    Odrv4 I__10410 (
            .O(N__45018),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    InMux I__10409 (
            .O(N__45015),
            .I(N__45012));
    LocalMux I__10408 (
            .O(N__45012),
            .I(N__45007));
    InMux I__10407 (
            .O(N__45011),
            .I(N__45004));
    InMux I__10406 (
            .O(N__45010),
            .I(N__45001));
    Span4Mux_h I__10405 (
            .O(N__45007),
            .I(N__44996));
    LocalMux I__10404 (
            .O(N__45004),
            .I(N__44996));
    LocalMux I__10403 (
            .O(N__45001),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    Odrv4 I__10402 (
            .O(N__44996),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    InMux I__10401 (
            .O(N__44991),
            .I(N__44987));
    InMux I__10400 (
            .O(N__44990),
            .I(N__44984));
    LocalMux I__10399 (
            .O(N__44987),
            .I(N__44980));
    LocalMux I__10398 (
            .O(N__44984),
            .I(N__44977));
    InMux I__10397 (
            .O(N__44983),
            .I(N__44973));
    Span4Mux_v I__10396 (
            .O(N__44980),
            .I(N__44968));
    Span4Mux_v I__10395 (
            .O(N__44977),
            .I(N__44968));
    InMux I__10394 (
            .O(N__44976),
            .I(N__44965));
    LocalMux I__10393 (
            .O(N__44973),
            .I(N__44962));
    Sp12to4 I__10392 (
            .O(N__44968),
            .I(N__44957));
    LocalMux I__10391 (
            .O(N__44965),
            .I(N__44957));
    Odrv4 I__10390 (
            .O(N__44962),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    Odrv12 I__10389 (
            .O(N__44957),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__10388 (
            .O(N__44952),
            .I(N__44949));
    LocalMux I__10387 (
            .O(N__44949),
            .I(N__44946));
    Span4Mux_h I__10386 (
            .O(N__44946),
            .I(N__44943));
    Odrv4 I__10385 (
            .O(N__44943),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    InMux I__10384 (
            .O(N__44940),
            .I(N__44937));
    LocalMux I__10383 (
            .O(N__44937),
            .I(N__44934));
    Odrv4 I__10382 (
            .O(N__44934),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt24 ));
    InMux I__10381 (
            .O(N__44931),
            .I(N__44926));
    InMux I__10380 (
            .O(N__44930),
            .I(N__44921));
    InMux I__10379 (
            .O(N__44929),
            .I(N__44921));
    LocalMux I__10378 (
            .O(N__44926),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    LocalMux I__10377 (
            .O(N__44921),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    CascadeMux I__10376 (
            .O(N__44916),
            .I(N__44911));
    InMux I__10375 (
            .O(N__44915),
            .I(N__44908));
    InMux I__10374 (
            .O(N__44914),
            .I(N__44903));
    InMux I__10373 (
            .O(N__44911),
            .I(N__44903));
    LocalMux I__10372 (
            .O(N__44908),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    LocalMux I__10371 (
            .O(N__44903),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    CascadeMux I__10370 (
            .O(N__44898),
            .I(N__44895));
    InMux I__10369 (
            .O(N__44895),
            .I(N__44892));
    LocalMux I__10368 (
            .O(N__44892),
            .I(N__44889));
    Odrv12 I__10367 (
            .O(N__44889),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ));
    InMux I__10366 (
            .O(N__44886),
            .I(N__44881));
    InMux I__10365 (
            .O(N__44885),
            .I(N__44878));
    InMux I__10364 (
            .O(N__44884),
            .I(N__44875));
    LocalMux I__10363 (
            .O(N__44881),
            .I(N__44872));
    LocalMux I__10362 (
            .O(N__44878),
            .I(N__44868));
    LocalMux I__10361 (
            .O(N__44875),
            .I(N__44865));
    Span4Mux_v I__10360 (
            .O(N__44872),
            .I(N__44862));
    InMux I__10359 (
            .O(N__44871),
            .I(N__44859));
    Span4Mux_v I__10358 (
            .O(N__44868),
            .I(N__44852));
    Span4Mux_v I__10357 (
            .O(N__44865),
            .I(N__44852));
    Span4Mux_h I__10356 (
            .O(N__44862),
            .I(N__44852));
    LocalMux I__10355 (
            .O(N__44859),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    Odrv4 I__10354 (
            .O(N__44852),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    CascadeMux I__10353 (
            .O(N__44847),
            .I(N__44844));
    InMux I__10352 (
            .O(N__44844),
            .I(N__44839));
    InMux I__10351 (
            .O(N__44843),
            .I(N__44834));
    InMux I__10350 (
            .O(N__44842),
            .I(N__44834));
    LocalMux I__10349 (
            .O(N__44839),
            .I(N__44831));
    LocalMux I__10348 (
            .O(N__44834),
            .I(N__44827));
    Span4Mux_v I__10347 (
            .O(N__44831),
            .I(N__44824));
    InMux I__10346 (
            .O(N__44830),
            .I(N__44821));
    Span4Mux_h I__10345 (
            .O(N__44827),
            .I(N__44818));
    Span4Mux_h I__10344 (
            .O(N__44824),
            .I(N__44815));
    LocalMux I__10343 (
            .O(N__44821),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__10342 (
            .O(N__44818),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__10341 (
            .O(N__44815),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__10340 (
            .O(N__44808),
            .I(N__44802));
    InMux I__10339 (
            .O(N__44807),
            .I(N__44799));
    InMux I__10338 (
            .O(N__44806),
            .I(N__44796));
    InMux I__10337 (
            .O(N__44805),
            .I(N__44793));
    LocalMux I__10336 (
            .O(N__44802),
            .I(N__44790));
    LocalMux I__10335 (
            .O(N__44799),
            .I(N__44787));
    LocalMux I__10334 (
            .O(N__44796),
            .I(N__44784));
    LocalMux I__10333 (
            .O(N__44793),
            .I(N__44779));
    Span12Mux_s6_v I__10332 (
            .O(N__44790),
            .I(N__44779));
    Span4Mux_v I__10331 (
            .O(N__44787),
            .I(N__44774));
    Span4Mux_h I__10330 (
            .O(N__44784),
            .I(N__44774));
    Odrv12 I__10329 (
            .O(N__44779),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__10328 (
            .O(N__44774),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__10327 (
            .O(N__44769),
            .I(N__44764));
    InMux I__10326 (
            .O(N__44768),
            .I(N__44761));
    InMux I__10325 (
            .O(N__44767),
            .I(N__44758));
    LocalMux I__10324 (
            .O(N__44764),
            .I(N__44755));
    LocalMux I__10323 (
            .O(N__44761),
            .I(N__44751));
    LocalMux I__10322 (
            .O(N__44758),
            .I(N__44746));
    Span4Mux_v I__10321 (
            .O(N__44755),
            .I(N__44746));
    InMux I__10320 (
            .O(N__44754),
            .I(N__44743));
    Span4Mux_h I__10319 (
            .O(N__44751),
            .I(N__44740));
    Sp12to4 I__10318 (
            .O(N__44746),
            .I(N__44735));
    LocalMux I__10317 (
            .O(N__44743),
            .I(N__44735));
    Odrv4 I__10316 (
            .O(N__44740),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv12 I__10315 (
            .O(N__44735),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    CascadeMux I__10314 (
            .O(N__44730),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ));
    InMux I__10313 (
            .O(N__44727),
            .I(N__44724));
    LocalMux I__10312 (
            .O(N__44724),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ));
    InMux I__10311 (
            .O(N__44721),
            .I(N__44718));
    LocalMux I__10310 (
            .O(N__44718),
            .I(N__44713));
    InMux I__10309 (
            .O(N__44717),
            .I(N__44710));
    InMux I__10308 (
            .O(N__44716),
            .I(N__44707));
    Span4Mux_v I__10307 (
            .O(N__44713),
            .I(N__44701));
    LocalMux I__10306 (
            .O(N__44710),
            .I(N__44701));
    LocalMux I__10305 (
            .O(N__44707),
            .I(N__44698));
    InMux I__10304 (
            .O(N__44706),
            .I(N__44695));
    Span4Mux_v I__10303 (
            .O(N__44701),
            .I(N__44692));
    Span4Mux_v I__10302 (
            .O(N__44698),
            .I(N__44689));
    LocalMux I__10301 (
            .O(N__44695),
            .I(N__44686));
    Span4Mux_h I__10300 (
            .O(N__44692),
            .I(N__44683));
    Odrv4 I__10299 (
            .O(N__44689),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv12 I__10298 (
            .O(N__44686),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__10297 (
            .O(N__44683),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__10296 (
            .O(N__44676),
            .I(N__44673));
    LocalMux I__10295 (
            .O(N__44673),
            .I(N__44670));
    Span4Mux_h I__10294 (
            .O(N__44670),
            .I(N__44667));
    Odrv4 I__10293 (
            .O(N__44667),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    CascadeMux I__10292 (
            .O(N__44664),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ));
    CascadeMux I__10291 (
            .O(N__44661),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__10290 (
            .O(N__44658),
            .I(N__44655));
    LocalMux I__10289 (
            .O(N__44655),
            .I(N__44652));
    Odrv4 I__10288 (
            .O(N__44652),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ));
    InMux I__10287 (
            .O(N__44649),
            .I(N__44646));
    LocalMux I__10286 (
            .O(N__44646),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ));
    InMux I__10285 (
            .O(N__44643),
            .I(N__44639));
    InMux I__10284 (
            .O(N__44642),
            .I(N__44635));
    LocalMux I__10283 (
            .O(N__44639),
            .I(N__44632));
    InMux I__10282 (
            .O(N__44638),
            .I(N__44629));
    LocalMux I__10281 (
            .O(N__44635),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    Odrv4 I__10280 (
            .O(N__44632),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    LocalMux I__10279 (
            .O(N__44629),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    InMux I__10278 (
            .O(N__44622),
            .I(N__44618));
    CascadeMux I__10277 (
            .O(N__44621),
            .I(N__44613));
    LocalMux I__10276 (
            .O(N__44618),
            .I(N__44610));
    InMux I__10275 (
            .O(N__44617),
            .I(N__44607));
    InMux I__10274 (
            .O(N__44616),
            .I(N__44604));
    InMux I__10273 (
            .O(N__44613),
            .I(N__44601));
    Span12Mux_h I__10272 (
            .O(N__44610),
            .I(N__44598));
    LocalMux I__10271 (
            .O(N__44607),
            .I(N__44591));
    LocalMux I__10270 (
            .O(N__44604),
            .I(N__44591));
    LocalMux I__10269 (
            .O(N__44601),
            .I(N__44591));
    Odrv12 I__10268 (
            .O(N__44598),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv12 I__10267 (
            .O(N__44591),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__10266 (
            .O(N__44586),
            .I(N__44583));
    LocalMux I__10265 (
            .O(N__44583),
            .I(N__44580));
    Span4Mux_h I__10264 (
            .O(N__44580),
            .I(N__44577));
    Odrv4 I__10263 (
            .O(N__44577),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__10262 (
            .O(N__44574),
            .I(N__44571));
    InMux I__10261 (
            .O(N__44571),
            .I(N__44567));
    InMux I__10260 (
            .O(N__44570),
            .I(N__44564));
    LocalMux I__10259 (
            .O(N__44567),
            .I(N__44558));
    LocalMux I__10258 (
            .O(N__44564),
            .I(N__44558));
    InMux I__10257 (
            .O(N__44563),
            .I(N__44555));
    Span4Mux_h I__10256 (
            .O(N__44558),
            .I(N__44552));
    LocalMux I__10255 (
            .O(N__44555),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__10254 (
            .O(N__44552),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__10253 (
            .O(N__44547),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__10252 (
            .O(N__44544),
            .I(N__44540));
    CascadeMux I__10251 (
            .O(N__44543),
            .I(N__44537));
    InMux I__10250 (
            .O(N__44540),
            .I(N__44531));
    InMux I__10249 (
            .O(N__44537),
            .I(N__44531));
    InMux I__10248 (
            .O(N__44536),
            .I(N__44528));
    LocalMux I__10247 (
            .O(N__44531),
            .I(N__44525));
    LocalMux I__10246 (
            .O(N__44528),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv12 I__10245 (
            .O(N__44525),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__10244 (
            .O(N__44520),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__10243 (
            .O(N__44517),
            .I(N__44513));
    InMux I__10242 (
            .O(N__44516),
            .I(N__44510));
    LocalMux I__10241 (
            .O(N__44513),
            .I(N__44507));
    LocalMux I__10240 (
            .O(N__44510),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv12 I__10239 (
            .O(N__44507),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__10238 (
            .O(N__44502),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__10237 (
            .O(N__44499),
            .I(N__44463));
    InMux I__10236 (
            .O(N__44498),
            .I(N__44463));
    InMux I__10235 (
            .O(N__44497),
            .I(N__44463));
    InMux I__10234 (
            .O(N__44496),
            .I(N__44454));
    InMux I__10233 (
            .O(N__44495),
            .I(N__44454));
    InMux I__10232 (
            .O(N__44494),
            .I(N__44454));
    InMux I__10231 (
            .O(N__44493),
            .I(N__44454));
    InMux I__10230 (
            .O(N__44492),
            .I(N__44445));
    InMux I__10229 (
            .O(N__44491),
            .I(N__44445));
    InMux I__10228 (
            .O(N__44490),
            .I(N__44445));
    InMux I__10227 (
            .O(N__44489),
            .I(N__44445));
    InMux I__10226 (
            .O(N__44488),
            .I(N__44436));
    InMux I__10225 (
            .O(N__44487),
            .I(N__44436));
    InMux I__10224 (
            .O(N__44486),
            .I(N__44436));
    InMux I__10223 (
            .O(N__44485),
            .I(N__44436));
    InMux I__10222 (
            .O(N__44484),
            .I(N__44427));
    InMux I__10221 (
            .O(N__44483),
            .I(N__44427));
    InMux I__10220 (
            .O(N__44482),
            .I(N__44427));
    InMux I__10219 (
            .O(N__44481),
            .I(N__44427));
    InMux I__10218 (
            .O(N__44480),
            .I(N__44420));
    InMux I__10217 (
            .O(N__44479),
            .I(N__44420));
    InMux I__10216 (
            .O(N__44478),
            .I(N__44420));
    InMux I__10215 (
            .O(N__44477),
            .I(N__44411));
    InMux I__10214 (
            .O(N__44476),
            .I(N__44411));
    InMux I__10213 (
            .O(N__44475),
            .I(N__44411));
    InMux I__10212 (
            .O(N__44474),
            .I(N__44411));
    InMux I__10211 (
            .O(N__44473),
            .I(N__44402));
    InMux I__10210 (
            .O(N__44472),
            .I(N__44402));
    InMux I__10209 (
            .O(N__44471),
            .I(N__44402));
    InMux I__10208 (
            .O(N__44470),
            .I(N__44402));
    LocalMux I__10207 (
            .O(N__44463),
            .I(N__44393));
    LocalMux I__10206 (
            .O(N__44454),
            .I(N__44393));
    LocalMux I__10205 (
            .O(N__44445),
            .I(N__44393));
    LocalMux I__10204 (
            .O(N__44436),
            .I(N__44393));
    LocalMux I__10203 (
            .O(N__44427),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__10202 (
            .O(N__44420),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__10201 (
            .O(N__44411),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__10200 (
            .O(N__44402),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__10199 (
            .O(N__44393),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__10198 (
            .O(N__44382),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__10197 (
            .O(N__44379),
            .I(N__44375));
    InMux I__10196 (
            .O(N__44378),
            .I(N__44372));
    LocalMux I__10195 (
            .O(N__44375),
            .I(N__44369));
    LocalMux I__10194 (
            .O(N__44372),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv12 I__10193 (
            .O(N__44369),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__10192 (
            .O(N__44364),
            .I(N__44360));
    CEMux I__10191 (
            .O(N__44363),
            .I(N__44357));
    LocalMux I__10190 (
            .O(N__44360),
            .I(N__44352));
    LocalMux I__10189 (
            .O(N__44357),
            .I(N__44349));
    CEMux I__10188 (
            .O(N__44356),
            .I(N__44346));
    CEMux I__10187 (
            .O(N__44355),
            .I(N__44343));
    Span4Mux_v I__10186 (
            .O(N__44352),
            .I(N__44338));
    Span4Mux_v I__10185 (
            .O(N__44349),
            .I(N__44338));
    LocalMux I__10184 (
            .O(N__44346),
            .I(N__44333));
    LocalMux I__10183 (
            .O(N__44343),
            .I(N__44333));
    Span4Mux_h I__10182 (
            .O(N__44338),
            .I(N__44328));
    Span4Mux_v I__10181 (
            .O(N__44333),
            .I(N__44328));
    Odrv4 I__10180 (
            .O(N__44328),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    InMux I__10179 (
            .O(N__44325),
            .I(N__44322));
    LocalMux I__10178 (
            .O(N__44322),
            .I(N__44317));
    InMux I__10177 (
            .O(N__44321),
            .I(N__44314));
    InMux I__10176 (
            .O(N__44320),
            .I(N__44311));
    Span4Mux_v I__10175 (
            .O(N__44317),
            .I(N__44308));
    LocalMux I__10174 (
            .O(N__44314),
            .I(N__44305));
    LocalMux I__10173 (
            .O(N__44311),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__10172 (
            .O(N__44308),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv12 I__10171 (
            .O(N__44305),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__10170 (
            .O(N__44298),
            .I(N__44293));
    InMux I__10169 (
            .O(N__44297),
            .I(N__44290));
    InMux I__10168 (
            .O(N__44296),
            .I(N__44287));
    LocalMux I__10167 (
            .O(N__44293),
            .I(N__44283));
    LocalMux I__10166 (
            .O(N__44290),
            .I(N__44278));
    LocalMux I__10165 (
            .O(N__44287),
            .I(N__44278));
    CascadeMux I__10164 (
            .O(N__44286),
            .I(N__44275));
    Span4Mux_h I__10163 (
            .O(N__44283),
            .I(N__44272));
    Span12Mux_h I__10162 (
            .O(N__44278),
            .I(N__44269));
    InMux I__10161 (
            .O(N__44275),
            .I(N__44266));
    Odrv4 I__10160 (
            .O(N__44272),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv12 I__10159 (
            .O(N__44269),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    LocalMux I__10158 (
            .O(N__44266),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__10157 (
            .O(N__44259),
            .I(N__44256));
    LocalMux I__10156 (
            .O(N__44256),
            .I(N__44252));
    InMux I__10155 (
            .O(N__44255),
            .I(N__44248));
    Span4Mux_h I__10154 (
            .O(N__44252),
            .I(N__44245));
    InMux I__10153 (
            .O(N__44251),
            .I(N__44242));
    LocalMux I__10152 (
            .O(N__44248),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__10151 (
            .O(N__44245),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    LocalMux I__10150 (
            .O(N__44242),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    InMux I__10149 (
            .O(N__44235),
            .I(N__44230));
    InMux I__10148 (
            .O(N__44234),
            .I(N__44227));
    InMux I__10147 (
            .O(N__44233),
            .I(N__44224));
    LocalMux I__10146 (
            .O(N__44230),
            .I(N__44221));
    LocalMux I__10145 (
            .O(N__44227),
            .I(N__44218));
    LocalMux I__10144 (
            .O(N__44224),
            .I(N__44213));
    Span4Mux_h I__10143 (
            .O(N__44221),
            .I(N__44213));
    Span4Mux_h I__10142 (
            .O(N__44218),
            .I(N__44210));
    Odrv4 I__10141 (
            .O(N__44213),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    Odrv4 I__10140 (
            .O(N__44210),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    InMux I__10139 (
            .O(N__44205),
            .I(N__44202));
    LocalMux I__10138 (
            .O(N__44202),
            .I(N__44197));
    InMux I__10137 (
            .O(N__44201),
            .I(N__44194));
    InMux I__10136 (
            .O(N__44200),
            .I(N__44191));
    Span4Mux_h I__10135 (
            .O(N__44197),
            .I(N__44188));
    LocalMux I__10134 (
            .O(N__44194),
            .I(N__44185));
    LocalMux I__10133 (
            .O(N__44191),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv4 I__10132 (
            .O(N__44188),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv12 I__10131 (
            .O(N__44185),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    CascadeMux I__10130 (
            .O(N__44178),
            .I(N__44175));
    InMux I__10129 (
            .O(N__44175),
            .I(N__44171));
    InMux I__10128 (
            .O(N__44174),
            .I(N__44168));
    LocalMux I__10127 (
            .O(N__44171),
            .I(N__44162));
    LocalMux I__10126 (
            .O(N__44168),
            .I(N__44162));
    InMux I__10125 (
            .O(N__44167),
            .I(N__44159));
    Span4Mux_h I__10124 (
            .O(N__44162),
            .I(N__44156));
    LocalMux I__10123 (
            .O(N__44159),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__10122 (
            .O(N__44156),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__10121 (
            .O(N__44151),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__10120 (
            .O(N__44148),
            .I(N__44144));
    CascadeMux I__10119 (
            .O(N__44147),
            .I(N__44141));
    InMux I__10118 (
            .O(N__44144),
            .I(N__44135));
    InMux I__10117 (
            .O(N__44141),
            .I(N__44135));
    InMux I__10116 (
            .O(N__44140),
            .I(N__44132));
    LocalMux I__10115 (
            .O(N__44135),
            .I(N__44129));
    LocalMux I__10114 (
            .O(N__44132),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv12 I__10113 (
            .O(N__44129),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__10112 (
            .O(N__44124),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__10111 (
            .O(N__44121),
            .I(N__44114));
    InMux I__10110 (
            .O(N__44120),
            .I(N__44114));
    InMux I__10109 (
            .O(N__44119),
            .I(N__44111));
    LocalMux I__10108 (
            .O(N__44114),
            .I(N__44108));
    LocalMux I__10107 (
            .O(N__44111),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv12 I__10106 (
            .O(N__44108),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__10105 (
            .O(N__44103),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__10104 (
            .O(N__44100),
            .I(N__44097));
    InMux I__10103 (
            .O(N__44097),
            .I(N__44092));
    InMux I__10102 (
            .O(N__44096),
            .I(N__44089));
    InMux I__10101 (
            .O(N__44095),
            .I(N__44086));
    LocalMux I__10100 (
            .O(N__44092),
            .I(N__44081));
    LocalMux I__10099 (
            .O(N__44089),
            .I(N__44081));
    LocalMux I__10098 (
            .O(N__44086),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv12 I__10097 (
            .O(N__44081),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__10096 (
            .O(N__44076),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__10095 (
            .O(N__44073),
            .I(N__44069));
    CascadeMux I__10094 (
            .O(N__44072),
            .I(N__44066));
    InMux I__10093 (
            .O(N__44069),
            .I(N__44060));
    InMux I__10092 (
            .O(N__44066),
            .I(N__44060));
    InMux I__10091 (
            .O(N__44065),
            .I(N__44057));
    LocalMux I__10090 (
            .O(N__44060),
            .I(N__44054));
    LocalMux I__10089 (
            .O(N__44057),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv12 I__10088 (
            .O(N__44054),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__10087 (
            .O(N__44049),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__10086 (
            .O(N__44046),
            .I(N__44039));
    InMux I__10085 (
            .O(N__44045),
            .I(N__44039));
    InMux I__10084 (
            .O(N__44044),
            .I(N__44036));
    LocalMux I__10083 (
            .O(N__44039),
            .I(N__44033));
    LocalMux I__10082 (
            .O(N__44036),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv12 I__10081 (
            .O(N__44033),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__10080 (
            .O(N__44028),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__10079 (
            .O(N__44025),
            .I(N__44022));
    InMux I__10078 (
            .O(N__44022),
            .I(N__44018));
    InMux I__10077 (
            .O(N__44021),
            .I(N__44015));
    LocalMux I__10076 (
            .O(N__44018),
            .I(N__44009));
    LocalMux I__10075 (
            .O(N__44015),
            .I(N__44009));
    InMux I__10074 (
            .O(N__44014),
            .I(N__44006));
    Span4Mux_v I__10073 (
            .O(N__44009),
            .I(N__44003));
    LocalMux I__10072 (
            .O(N__44006),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__10071 (
            .O(N__44003),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__10070 (
            .O(N__43998),
            .I(bfn_17_22_0_));
    InMux I__10069 (
            .O(N__43995),
            .I(N__43991));
    CascadeMux I__10068 (
            .O(N__43994),
            .I(N__43988));
    LocalMux I__10067 (
            .O(N__43991),
            .I(N__43984));
    InMux I__10066 (
            .O(N__43988),
            .I(N__43981));
    InMux I__10065 (
            .O(N__43987),
            .I(N__43978));
    Span4Mux_h I__10064 (
            .O(N__43984),
            .I(N__43975));
    LocalMux I__10063 (
            .O(N__43981),
            .I(N__43972));
    LocalMux I__10062 (
            .O(N__43978),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__10061 (
            .O(N__43975),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv12 I__10060 (
            .O(N__43972),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__10059 (
            .O(N__43965),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__10058 (
            .O(N__43962),
            .I(N__43959));
    InMux I__10057 (
            .O(N__43959),
            .I(N__43956));
    LocalMux I__10056 (
            .O(N__43956),
            .I(N__43951));
    InMux I__10055 (
            .O(N__43955),
            .I(N__43948));
    InMux I__10054 (
            .O(N__43954),
            .I(N__43945));
    Span4Mux_h I__10053 (
            .O(N__43951),
            .I(N__43942));
    LocalMux I__10052 (
            .O(N__43948),
            .I(N__43939));
    LocalMux I__10051 (
            .O(N__43945),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__10050 (
            .O(N__43942),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv12 I__10049 (
            .O(N__43939),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__10048 (
            .O(N__43932),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__10047 (
            .O(N__43929),
            .I(N__43922));
    InMux I__10046 (
            .O(N__43928),
            .I(N__43922));
    InMux I__10045 (
            .O(N__43927),
            .I(N__43919));
    LocalMux I__10044 (
            .O(N__43922),
            .I(N__43916));
    LocalMux I__10043 (
            .O(N__43919),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv12 I__10042 (
            .O(N__43916),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__10041 (
            .O(N__43911),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__10040 (
            .O(N__43908),
            .I(N__43902));
    InMux I__10039 (
            .O(N__43907),
            .I(N__43902));
    LocalMux I__10038 (
            .O(N__43902),
            .I(N__43898));
    InMux I__10037 (
            .O(N__43901),
            .I(N__43895));
    Span4Mux_h I__10036 (
            .O(N__43898),
            .I(N__43892));
    LocalMux I__10035 (
            .O(N__43895),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__10034 (
            .O(N__43892),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__10033 (
            .O(N__43887),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__10032 (
            .O(N__43884),
            .I(N__43880));
    InMux I__10031 (
            .O(N__43883),
            .I(N__43876));
    InMux I__10030 (
            .O(N__43880),
            .I(N__43873));
    InMux I__10029 (
            .O(N__43879),
            .I(N__43870));
    LocalMux I__10028 (
            .O(N__43876),
            .I(N__43865));
    LocalMux I__10027 (
            .O(N__43873),
            .I(N__43865));
    LocalMux I__10026 (
            .O(N__43870),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv12 I__10025 (
            .O(N__43865),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__10024 (
            .O(N__43860),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__10023 (
            .O(N__43857),
            .I(N__43853));
    CascadeMux I__10022 (
            .O(N__43856),
            .I(N__43850));
    InMux I__10021 (
            .O(N__43853),
            .I(N__43845));
    InMux I__10020 (
            .O(N__43850),
            .I(N__43845));
    LocalMux I__10019 (
            .O(N__43845),
            .I(N__43841));
    InMux I__10018 (
            .O(N__43844),
            .I(N__43838));
    Span4Mux_h I__10017 (
            .O(N__43841),
            .I(N__43835));
    LocalMux I__10016 (
            .O(N__43838),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__10015 (
            .O(N__43835),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__10014 (
            .O(N__43830),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__10013 (
            .O(N__43827),
            .I(N__43823));
    CascadeMux I__10012 (
            .O(N__43826),
            .I(N__43820));
    InMux I__10011 (
            .O(N__43823),
            .I(N__43815));
    InMux I__10010 (
            .O(N__43820),
            .I(N__43815));
    LocalMux I__10009 (
            .O(N__43815),
            .I(N__43811));
    InMux I__10008 (
            .O(N__43814),
            .I(N__43808));
    Span4Mux_v I__10007 (
            .O(N__43811),
            .I(N__43805));
    LocalMux I__10006 (
            .O(N__43808),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__10005 (
            .O(N__43805),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__10004 (
            .O(N__43800),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__10003 (
            .O(N__43797),
            .I(N__43791));
    InMux I__10002 (
            .O(N__43796),
            .I(N__43791));
    LocalMux I__10001 (
            .O(N__43791),
            .I(N__43787));
    InMux I__10000 (
            .O(N__43790),
            .I(N__43784));
    Span4Mux_v I__9999 (
            .O(N__43787),
            .I(N__43781));
    LocalMux I__9998 (
            .O(N__43784),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__9997 (
            .O(N__43781),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__9996 (
            .O(N__43776),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__9995 (
            .O(N__43773),
            .I(N__43770));
    InMux I__9994 (
            .O(N__43770),
            .I(N__43766));
    InMux I__9993 (
            .O(N__43769),
            .I(N__43763));
    LocalMux I__9992 (
            .O(N__43766),
            .I(N__43757));
    LocalMux I__9991 (
            .O(N__43763),
            .I(N__43757));
    InMux I__9990 (
            .O(N__43762),
            .I(N__43754));
    Span4Mux_v I__9989 (
            .O(N__43757),
            .I(N__43751));
    LocalMux I__9988 (
            .O(N__43754),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__9987 (
            .O(N__43751),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__9986 (
            .O(N__43746),
            .I(bfn_17_21_0_));
    CascadeMux I__9985 (
            .O(N__43743),
            .I(N__43739));
    InMux I__9984 (
            .O(N__43742),
            .I(N__43736));
    InMux I__9983 (
            .O(N__43739),
            .I(N__43733));
    LocalMux I__9982 (
            .O(N__43736),
            .I(N__43729));
    LocalMux I__9981 (
            .O(N__43733),
            .I(N__43726));
    InMux I__9980 (
            .O(N__43732),
            .I(N__43723));
    Span4Mux_v I__9979 (
            .O(N__43729),
            .I(N__43718));
    Span4Mux_v I__9978 (
            .O(N__43726),
            .I(N__43718));
    LocalMux I__9977 (
            .O(N__43723),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__9976 (
            .O(N__43718),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__9975 (
            .O(N__43713),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__9974 (
            .O(N__43710),
            .I(N__43707));
    LocalMux I__9973 (
            .O(N__43707),
            .I(N__43703));
    InMux I__9972 (
            .O(N__43706),
            .I(N__43699));
    Span4Mux_h I__9971 (
            .O(N__43703),
            .I(N__43696));
    InMux I__9970 (
            .O(N__43702),
            .I(N__43693));
    LocalMux I__9969 (
            .O(N__43699),
            .I(N__43690));
    Odrv4 I__9968 (
            .O(N__43696),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__9967 (
            .O(N__43693),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv12 I__9966 (
            .O(N__43690),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__9965 (
            .O(N__43683),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__9964 (
            .O(N__43680),
            .I(N__43676));
    CascadeMux I__9963 (
            .O(N__43679),
            .I(N__43673));
    LocalMux I__9962 (
            .O(N__43676),
            .I(N__43669));
    InMux I__9961 (
            .O(N__43673),
            .I(N__43666));
    InMux I__9960 (
            .O(N__43672),
            .I(N__43663));
    Sp12to4 I__9959 (
            .O(N__43669),
            .I(N__43658));
    LocalMux I__9958 (
            .O(N__43666),
            .I(N__43658));
    LocalMux I__9957 (
            .O(N__43663),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__9956 (
            .O(N__43658),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__9955 (
            .O(N__43653),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    CascadeMux I__9954 (
            .O(N__43650),
            .I(N__43646));
    InMux I__9953 (
            .O(N__43649),
            .I(N__43643));
    InMux I__9952 (
            .O(N__43646),
            .I(N__43640));
    LocalMux I__9951 (
            .O(N__43643),
            .I(N__43634));
    LocalMux I__9950 (
            .O(N__43640),
            .I(N__43634));
    InMux I__9949 (
            .O(N__43639),
            .I(N__43631));
    Span4Mux_v I__9948 (
            .O(N__43634),
            .I(N__43628));
    LocalMux I__9947 (
            .O(N__43631),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__9946 (
            .O(N__43628),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__9945 (
            .O(N__43623),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__9944 (
            .O(N__43620),
            .I(N__43616));
    CascadeMux I__9943 (
            .O(N__43619),
            .I(N__43613));
    InMux I__9942 (
            .O(N__43616),
            .I(N__43608));
    InMux I__9941 (
            .O(N__43613),
            .I(N__43608));
    LocalMux I__9940 (
            .O(N__43608),
            .I(N__43604));
    InMux I__9939 (
            .O(N__43607),
            .I(N__43601));
    Span4Mux_v I__9938 (
            .O(N__43604),
            .I(N__43598));
    LocalMux I__9937 (
            .O(N__43601),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__9936 (
            .O(N__43598),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__9935 (
            .O(N__43593),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__9934 (
            .O(N__43590),
            .I(N__43586));
    CascadeMux I__9933 (
            .O(N__43589),
            .I(N__43583));
    InMux I__9932 (
            .O(N__43586),
            .I(N__43578));
    InMux I__9931 (
            .O(N__43583),
            .I(N__43578));
    LocalMux I__9930 (
            .O(N__43578),
            .I(N__43574));
    InMux I__9929 (
            .O(N__43577),
            .I(N__43571));
    Span4Mux_h I__9928 (
            .O(N__43574),
            .I(N__43568));
    LocalMux I__9927 (
            .O(N__43571),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__9926 (
            .O(N__43568),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__9925 (
            .O(N__43563),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__9924 (
            .O(N__43560),
            .I(N__43554));
    InMux I__9923 (
            .O(N__43559),
            .I(N__43554));
    LocalMux I__9922 (
            .O(N__43554),
            .I(N__43550));
    InMux I__9921 (
            .O(N__43553),
            .I(N__43547));
    Span4Mux_v I__9920 (
            .O(N__43550),
            .I(N__43544));
    LocalMux I__9919 (
            .O(N__43547),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__9918 (
            .O(N__43544),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__9917 (
            .O(N__43539),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    CascadeMux I__9916 (
            .O(N__43536),
            .I(N__43533));
    InMux I__9915 (
            .O(N__43533),
            .I(N__43529));
    InMux I__9914 (
            .O(N__43532),
            .I(N__43526));
    LocalMux I__9913 (
            .O(N__43529),
            .I(N__43520));
    LocalMux I__9912 (
            .O(N__43526),
            .I(N__43520));
    InMux I__9911 (
            .O(N__43525),
            .I(N__43517));
    Span4Mux_v I__9910 (
            .O(N__43520),
            .I(N__43514));
    LocalMux I__9909 (
            .O(N__43517),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__9908 (
            .O(N__43514),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__9907 (
            .O(N__43509),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__9906 (
            .O(N__43506),
            .I(N__43502));
    CascadeMux I__9905 (
            .O(N__43505),
            .I(N__43499));
    InMux I__9904 (
            .O(N__43502),
            .I(N__43496));
    InMux I__9903 (
            .O(N__43499),
            .I(N__43493));
    LocalMux I__9902 (
            .O(N__43496),
            .I(N__43487));
    LocalMux I__9901 (
            .O(N__43493),
            .I(N__43487));
    InMux I__9900 (
            .O(N__43492),
            .I(N__43484));
    Span4Mux_v I__9899 (
            .O(N__43487),
            .I(N__43481));
    LocalMux I__9898 (
            .O(N__43484),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__9897 (
            .O(N__43481),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__9896 (
            .O(N__43476),
            .I(bfn_17_20_0_));
    InMux I__9895 (
            .O(N__43473),
            .I(N__43468));
    InMux I__9894 (
            .O(N__43472),
            .I(N__43465));
    InMux I__9893 (
            .O(N__43471),
            .I(N__43462));
    LocalMux I__9892 (
            .O(N__43468),
            .I(N__43459));
    LocalMux I__9891 (
            .O(N__43465),
            .I(N__43456));
    LocalMux I__9890 (
            .O(N__43462),
            .I(N__43453));
    Span4Mux_h I__9889 (
            .O(N__43459),
            .I(N__43449));
    Span4Mux_h I__9888 (
            .O(N__43456),
            .I(N__43446));
    Span4Mux_h I__9887 (
            .O(N__43453),
            .I(N__43443));
    InMux I__9886 (
            .O(N__43452),
            .I(N__43440));
    Odrv4 I__9885 (
            .O(N__43449),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__9884 (
            .O(N__43446),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__9883 (
            .O(N__43443),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__9882 (
            .O(N__43440),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__9881 (
            .O(N__43431),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__9880 (
            .O(N__43428),
            .I(N__43423));
    InMux I__9879 (
            .O(N__43427),
            .I(N__43420));
    InMux I__9878 (
            .O(N__43426),
            .I(N__43417));
    LocalMux I__9877 (
            .O(N__43423),
            .I(N__43413));
    LocalMux I__9876 (
            .O(N__43420),
            .I(N__43408));
    LocalMux I__9875 (
            .O(N__43417),
            .I(N__43408));
    InMux I__9874 (
            .O(N__43416),
            .I(N__43405));
    Span4Mux_v I__9873 (
            .O(N__43413),
            .I(N__43398));
    Span4Mux_v I__9872 (
            .O(N__43408),
            .I(N__43398));
    LocalMux I__9871 (
            .O(N__43405),
            .I(N__43398));
    Odrv4 I__9870 (
            .O(N__43398),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__9869 (
            .O(N__43395),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__9868 (
            .O(N__43392),
            .I(N__43387));
    InMux I__9867 (
            .O(N__43391),
            .I(N__43384));
    InMux I__9866 (
            .O(N__43390),
            .I(N__43381));
    LocalMux I__9865 (
            .O(N__43387),
            .I(N__43376));
    LocalMux I__9864 (
            .O(N__43384),
            .I(N__43376));
    LocalMux I__9863 (
            .O(N__43381),
            .I(N__43373));
    Span4Mux_v I__9862 (
            .O(N__43376),
            .I(N__43369));
    Span4Mux_h I__9861 (
            .O(N__43373),
            .I(N__43366));
    InMux I__9860 (
            .O(N__43372),
            .I(N__43363));
    Odrv4 I__9859 (
            .O(N__43369),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__9858 (
            .O(N__43366),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__9857 (
            .O(N__43363),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__9856 (
            .O(N__43356),
            .I(bfn_17_18_0_));
    InMux I__9855 (
            .O(N__43353),
            .I(N__43347));
    InMux I__9854 (
            .O(N__43352),
            .I(N__43347));
    LocalMux I__9853 (
            .O(N__43347),
            .I(N__43343));
    InMux I__9852 (
            .O(N__43346),
            .I(N__43340));
    Span4Mux_v I__9851 (
            .O(N__43343),
            .I(N__43335));
    LocalMux I__9850 (
            .O(N__43340),
            .I(N__43335));
    Span4Mux_h I__9849 (
            .O(N__43335),
            .I(N__43331));
    InMux I__9848 (
            .O(N__43334),
            .I(N__43328));
    Odrv4 I__9847 (
            .O(N__43331),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__9846 (
            .O(N__43328),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__9845 (
            .O(N__43323),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__9844 (
            .O(N__43320),
            .I(N__43316));
    InMux I__9843 (
            .O(N__43319),
            .I(N__43313));
    LocalMux I__9842 (
            .O(N__43316),
            .I(N__43307));
    LocalMux I__9841 (
            .O(N__43313),
            .I(N__43307));
    InMux I__9840 (
            .O(N__43312),
            .I(N__43304));
    Span4Mux_v I__9839 (
            .O(N__43307),
            .I(N__43298));
    LocalMux I__9838 (
            .O(N__43304),
            .I(N__43298));
    InMux I__9837 (
            .O(N__43303),
            .I(N__43295));
    Span4Mux_h I__9836 (
            .O(N__43298),
            .I(N__43292));
    LocalMux I__9835 (
            .O(N__43295),
            .I(N__43289));
    Odrv4 I__9834 (
            .O(N__43292),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv12 I__9833 (
            .O(N__43289),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__9832 (
            .O(N__43284),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__9831 (
            .O(N__43281),
            .I(N__43277));
    CascadeMux I__9830 (
            .O(N__43280),
            .I(N__43274));
    LocalMux I__9829 (
            .O(N__43277),
            .I(N__43270));
    InMux I__9828 (
            .O(N__43274),
            .I(N__43267));
    InMux I__9827 (
            .O(N__43273),
            .I(N__43264));
    Span4Mux_v I__9826 (
            .O(N__43270),
            .I(N__43261));
    LocalMux I__9825 (
            .O(N__43267),
            .I(N__43258));
    LocalMux I__9824 (
            .O(N__43264),
            .I(N__43255));
    Span4Mux_h I__9823 (
            .O(N__43261),
            .I(N__43249));
    Span4Mux_v I__9822 (
            .O(N__43258),
            .I(N__43249));
    Span4Mux_h I__9821 (
            .O(N__43255),
            .I(N__43246));
    InMux I__9820 (
            .O(N__43254),
            .I(N__43243));
    Odrv4 I__9819 (
            .O(N__43249),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__9818 (
            .O(N__43246),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__9817 (
            .O(N__43243),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__9816 (
            .O(N__43236),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    CEMux I__9815 (
            .O(N__43233),
            .I(N__43209));
    CEMux I__9814 (
            .O(N__43232),
            .I(N__43209));
    CEMux I__9813 (
            .O(N__43231),
            .I(N__43209));
    CEMux I__9812 (
            .O(N__43230),
            .I(N__43209));
    CEMux I__9811 (
            .O(N__43229),
            .I(N__43209));
    CEMux I__9810 (
            .O(N__43228),
            .I(N__43209));
    CEMux I__9809 (
            .O(N__43227),
            .I(N__43209));
    CEMux I__9808 (
            .O(N__43226),
            .I(N__43209));
    GlobalMux I__9807 (
            .O(N__43209),
            .I(N__43206));
    gio2CtrlBuf I__9806 (
            .O(N__43206),
            .I(\current_shift_inst.timer_s1.N_162_i_g ));
    InMux I__9805 (
            .O(N__43203),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__9804 (
            .O(N__43200),
            .I(N__43197));
    LocalMux I__9803 (
            .O(N__43197),
            .I(N__43194));
    Span4Mux_v I__9802 (
            .O(N__43194),
            .I(N__43189));
    InMux I__9801 (
            .O(N__43193),
            .I(N__43186));
    InMux I__9800 (
            .O(N__43192),
            .I(N__43183));
    Span4Mux_v I__9799 (
            .O(N__43189),
            .I(N__43176));
    LocalMux I__9798 (
            .O(N__43186),
            .I(N__43176));
    LocalMux I__9797 (
            .O(N__43183),
            .I(N__43176));
    Span4Mux_v I__9796 (
            .O(N__43176),
            .I(N__43173));
    Odrv4 I__9795 (
            .O(N__43173),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__9794 (
            .O(N__43170),
            .I(N__43167));
    LocalMux I__9793 (
            .O(N__43167),
            .I(N__43163));
    InMux I__9792 (
            .O(N__43166),
            .I(N__43159));
    Span12Mux_v I__9791 (
            .O(N__43163),
            .I(N__43156));
    InMux I__9790 (
            .O(N__43162),
            .I(N__43153));
    LocalMux I__9789 (
            .O(N__43159),
            .I(N__43150));
    Odrv12 I__9788 (
            .O(N__43156),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__9787 (
            .O(N__43153),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv12 I__9786 (
            .O(N__43150),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__9785 (
            .O(N__43143),
            .I(bfn_17_19_0_));
    CascadeMux I__9784 (
            .O(N__43140),
            .I(N__43136));
    InMux I__9783 (
            .O(N__43139),
            .I(N__43133));
    InMux I__9782 (
            .O(N__43136),
            .I(N__43129));
    LocalMux I__9781 (
            .O(N__43133),
            .I(N__43126));
    InMux I__9780 (
            .O(N__43132),
            .I(N__43123));
    LocalMux I__9779 (
            .O(N__43129),
            .I(N__43120));
    Span4Mux_h I__9778 (
            .O(N__43126),
            .I(N__43115));
    LocalMux I__9777 (
            .O(N__43123),
            .I(N__43115));
    Span4Mux_h I__9776 (
            .O(N__43120),
            .I(N__43111));
    Span4Mux_v I__9775 (
            .O(N__43115),
            .I(N__43108));
    InMux I__9774 (
            .O(N__43114),
            .I(N__43105));
    Odrv4 I__9773 (
            .O(N__43111),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__9772 (
            .O(N__43108),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__9771 (
            .O(N__43105),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__9770 (
            .O(N__43098),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__9769 (
            .O(N__43095),
            .I(N__43092));
    InMux I__9768 (
            .O(N__43092),
            .I(N__43089));
    LocalMux I__9767 (
            .O(N__43089),
            .I(N__43084));
    InMux I__9766 (
            .O(N__43088),
            .I(N__43081));
    InMux I__9765 (
            .O(N__43087),
            .I(N__43078));
    Span4Mux_v I__9764 (
            .O(N__43084),
            .I(N__43075));
    LocalMux I__9763 (
            .O(N__43081),
            .I(N__43070));
    LocalMux I__9762 (
            .O(N__43078),
            .I(N__43070));
    Span4Mux_h I__9761 (
            .O(N__43075),
            .I(N__43066));
    Span4Mux_h I__9760 (
            .O(N__43070),
            .I(N__43063));
    InMux I__9759 (
            .O(N__43069),
            .I(N__43060));
    Odrv4 I__9758 (
            .O(N__43066),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__9757 (
            .O(N__43063),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__9756 (
            .O(N__43060),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__9755 (
            .O(N__43053),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__9754 (
            .O(N__43050),
            .I(N__43047));
    InMux I__9753 (
            .O(N__43047),
            .I(N__43043));
    InMux I__9752 (
            .O(N__43046),
            .I(N__43039));
    LocalMux I__9751 (
            .O(N__43043),
            .I(N__43036));
    InMux I__9750 (
            .O(N__43042),
            .I(N__43033));
    LocalMux I__9749 (
            .O(N__43039),
            .I(N__43030));
    Span4Mux_v I__9748 (
            .O(N__43036),
            .I(N__43024));
    LocalMux I__9747 (
            .O(N__43033),
            .I(N__43024));
    Span4Mux_h I__9746 (
            .O(N__43030),
            .I(N__43021));
    InMux I__9745 (
            .O(N__43029),
            .I(N__43018));
    Odrv4 I__9744 (
            .O(N__43024),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__9743 (
            .O(N__43021),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__9742 (
            .O(N__43018),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__9741 (
            .O(N__43011),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__9740 (
            .O(N__43008),
            .I(N__43004));
    InMux I__9739 (
            .O(N__43007),
            .I(N__43001));
    InMux I__9738 (
            .O(N__43004),
            .I(N__42998));
    LocalMux I__9737 (
            .O(N__43001),
            .I(N__42994));
    LocalMux I__9736 (
            .O(N__42998),
            .I(N__42991));
    InMux I__9735 (
            .O(N__42997),
            .I(N__42988));
    Span4Mux_h I__9734 (
            .O(N__42994),
            .I(N__42981));
    Span4Mux_v I__9733 (
            .O(N__42991),
            .I(N__42981));
    LocalMux I__9732 (
            .O(N__42988),
            .I(N__42981));
    Span4Mux_h I__9731 (
            .O(N__42981),
            .I(N__42977));
    InMux I__9730 (
            .O(N__42980),
            .I(N__42974));
    Odrv4 I__9729 (
            .O(N__42977),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__9728 (
            .O(N__42974),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__9727 (
            .O(N__42969),
            .I(bfn_17_17_0_));
    InMux I__9726 (
            .O(N__42966),
            .I(N__42960));
    InMux I__9725 (
            .O(N__42965),
            .I(N__42960));
    LocalMux I__9724 (
            .O(N__42960),
            .I(N__42956));
    InMux I__9723 (
            .O(N__42959),
            .I(N__42953));
    Span4Mux_v I__9722 (
            .O(N__42956),
            .I(N__42948));
    LocalMux I__9721 (
            .O(N__42953),
            .I(N__42948));
    Span4Mux_h I__9720 (
            .O(N__42948),
            .I(N__42944));
    InMux I__9719 (
            .O(N__42947),
            .I(N__42941));
    Odrv4 I__9718 (
            .O(N__42944),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__9717 (
            .O(N__42941),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__9716 (
            .O(N__42936),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__9715 (
            .O(N__42933),
            .I(N__42928));
    InMux I__9714 (
            .O(N__42932),
            .I(N__42925));
    InMux I__9713 (
            .O(N__42931),
            .I(N__42922));
    LocalMux I__9712 (
            .O(N__42928),
            .I(N__42917));
    LocalMux I__9711 (
            .O(N__42925),
            .I(N__42917));
    LocalMux I__9710 (
            .O(N__42922),
            .I(N__42914));
    Span4Mux_h I__9709 (
            .O(N__42917),
            .I(N__42910));
    Span4Mux_h I__9708 (
            .O(N__42914),
            .I(N__42907));
    InMux I__9707 (
            .O(N__42913),
            .I(N__42904));
    Odrv4 I__9706 (
            .O(N__42910),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__9705 (
            .O(N__42907),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__9704 (
            .O(N__42904),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__9703 (
            .O(N__42897),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__9702 (
            .O(N__42894),
            .I(N__42889));
    InMux I__9701 (
            .O(N__42893),
            .I(N__42886));
    InMux I__9700 (
            .O(N__42892),
            .I(N__42883));
    LocalMux I__9699 (
            .O(N__42889),
            .I(N__42880));
    LocalMux I__9698 (
            .O(N__42886),
            .I(N__42875));
    LocalMux I__9697 (
            .O(N__42883),
            .I(N__42875));
    Span4Mux_v I__9696 (
            .O(N__42880),
            .I(N__42869));
    Span4Mux_v I__9695 (
            .O(N__42875),
            .I(N__42869));
    InMux I__9694 (
            .O(N__42874),
            .I(N__42866));
    Odrv4 I__9693 (
            .O(N__42869),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__9692 (
            .O(N__42866),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__9691 (
            .O(N__42861),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__9690 (
            .O(N__42858),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__9689 (
            .O(N__42855),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__9688 (
            .O(N__42852),
            .I(N__42848));
    CascadeMux I__9687 (
            .O(N__42851),
            .I(N__42845));
    InMux I__9686 (
            .O(N__42848),
            .I(N__42842));
    InMux I__9685 (
            .O(N__42845),
            .I(N__42839));
    LocalMux I__9684 (
            .O(N__42842),
            .I(N__42835));
    LocalMux I__9683 (
            .O(N__42839),
            .I(N__42832));
    InMux I__9682 (
            .O(N__42838),
            .I(N__42829));
    Span4Mux_v I__9681 (
            .O(N__42835),
            .I(N__42826));
    Span4Mux_v I__9680 (
            .O(N__42832),
            .I(N__42821));
    LocalMux I__9679 (
            .O(N__42829),
            .I(N__42821));
    Span4Mux_h I__9678 (
            .O(N__42826),
            .I(N__42817));
    Span4Mux_h I__9677 (
            .O(N__42821),
            .I(N__42814));
    InMux I__9676 (
            .O(N__42820),
            .I(N__42811));
    Odrv4 I__9675 (
            .O(N__42817),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__9674 (
            .O(N__42814),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__9673 (
            .O(N__42811),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__9672 (
            .O(N__42804),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__9671 (
            .O(N__42801),
            .I(N__42797));
    InMux I__9670 (
            .O(N__42800),
            .I(N__42793));
    InMux I__9669 (
            .O(N__42797),
            .I(N__42790));
    InMux I__9668 (
            .O(N__42796),
            .I(N__42787));
    LocalMux I__9667 (
            .O(N__42793),
            .I(N__42784));
    LocalMux I__9666 (
            .O(N__42790),
            .I(N__42781));
    LocalMux I__9665 (
            .O(N__42787),
            .I(N__42778));
    Span4Mux_h I__9664 (
            .O(N__42784),
            .I(N__42774));
    Span4Mux_v I__9663 (
            .O(N__42781),
            .I(N__42769));
    Span4Mux_v I__9662 (
            .O(N__42778),
            .I(N__42769));
    InMux I__9661 (
            .O(N__42777),
            .I(N__42766));
    Odrv4 I__9660 (
            .O(N__42774),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__9659 (
            .O(N__42769),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__9658 (
            .O(N__42766),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__9657 (
            .O(N__42759),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__9656 (
            .O(N__42756),
            .I(N__42752));
    InMux I__9655 (
            .O(N__42755),
            .I(N__42749));
    InMux I__9654 (
            .O(N__42752),
            .I(N__42746));
    LocalMux I__9653 (
            .O(N__42749),
            .I(N__42743));
    LocalMux I__9652 (
            .O(N__42746),
            .I(N__42739));
    Span4Mux_v I__9651 (
            .O(N__42743),
            .I(N__42736));
    InMux I__9650 (
            .O(N__42742),
            .I(N__42733));
    Span4Mux_v I__9649 (
            .O(N__42739),
            .I(N__42725));
    Span4Mux_h I__9648 (
            .O(N__42736),
            .I(N__42725));
    LocalMux I__9647 (
            .O(N__42733),
            .I(N__42725));
    InMux I__9646 (
            .O(N__42732),
            .I(N__42722));
    Odrv4 I__9645 (
            .O(N__42725),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__9644 (
            .O(N__42722),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__9643 (
            .O(N__42717),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__9642 (
            .O(N__42714),
            .I(N__42711));
    InMux I__9641 (
            .O(N__42711),
            .I(N__42706));
    InMux I__9640 (
            .O(N__42710),
            .I(N__42701));
    InMux I__9639 (
            .O(N__42709),
            .I(N__42701));
    LocalMux I__9638 (
            .O(N__42706),
            .I(N__42698));
    LocalMux I__9637 (
            .O(N__42701),
            .I(N__42695));
    Span12Mux_v I__9636 (
            .O(N__42698),
            .I(N__42691));
    Span4Mux_v I__9635 (
            .O(N__42695),
            .I(N__42688));
    InMux I__9634 (
            .O(N__42694),
            .I(N__42685));
    Odrv12 I__9633 (
            .O(N__42691),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__9632 (
            .O(N__42688),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__9631 (
            .O(N__42685),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__9630 (
            .O(N__42678),
            .I(bfn_17_16_0_));
    InMux I__9629 (
            .O(N__42675),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__9628 (
            .O(N__42672),
            .I(N__42667));
    InMux I__9627 (
            .O(N__42671),
            .I(N__42664));
    InMux I__9626 (
            .O(N__42670),
            .I(N__42661));
    InMux I__9625 (
            .O(N__42667),
            .I(N__42658));
    LocalMux I__9624 (
            .O(N__42664),
            .I(N__42655));
    LocalMux I__9623 (
            .O(N__42661),
            .I(N__42652));
    LocalMux I__9622 (
            .O(N__42658),
            .I(N__42648));
    Span4Mux_v I__9621 (
            .O(N__42655),
            .I(N__42643));
    Span4Mux_v I__9620 (
            .O(N__42652),
            .I(N__42643));
    InMux I__9619 (
            .O(N__42651),
            .I(N__42640));
    Span12Mux_v I__9618 (
            .O(N__42648),
            .I(N__42637));
    Span4Mux_h I__9617 (
            .O(N__42643),
            .I(N__42634));
    LocalMux I__9616 (
            .O(N__42640),
            .I(N__42631));
    Odrv12 I__9615 (
            .O(N__42637),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__9614 (
            .O(N__42634),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__9613 (
            .O(N__42631),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__9612 (
            .O(N__42624),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__9611 (
            .O(N__42621),
            .I(N__42617));
    InMux I__9610 (
            .O(N__42620),
            .I(N__42614));
    LocalMux I__9609 (
            .O(N__42617),
            .I(N__42608));
    LocalMux I__9608 (
            .O(N__42614),
            .I(N__42608));
    InMux I__9607 (
            .O(N__42613),
            .I(N__42605));
    Span4Mux_v I__9606 (
            .O(N__42608),
            .I(N__42599));
    LocalMux I__9605 (
            .O(N__42605),
            .I(N__42599));
    InMux I__9604 (
            .O(N__42604),
            .I(N__42596));
    Span4Mux_h I__9603 (
            .O(N__42599),
            .I(N__42593));
    LocalMux I__9602 (
            .O(N__42596),
            .I(N__42590));
    Odrv4 I__9601 (
            .O(N__42593),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__9600 (
            .O(N__42590),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__9599 (
            .O(N__42585),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__9598 (
            .O(N__42582),
            .I(N__42578));
    InMux I__9597 (
            .O(N__42581),
            .I(N__42573));
    InMux I__9596 (
            .O(N__42578),
            .I(N__42568));
    InMux I__9595 (
            .O(N__42577),
            .I(N__42568));
    InMux I__9594 (
            .O(N__42576),
            .I(N__42565));
    LocalMux I__9593 (
            .O(N__42573),
            .I(N__42562));
    LocalMux I__9592 (
            .O(N__42568),
            .I(N__42557));
    LocalMux I__9591 (
            .O(N__42565),
            .I(N__42557));
    Span4Mux_v I__9590 (
            .O(N__42562),
            .I(N__42554));
    Span4Mux_v I__9589 (
            .O(N__42557),
            .I(N__42551));
    Odrv4 I__9588 (
            .O(N__42554),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__9587 (
            .O(N__42551),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__9586 (
            .O(N__42546),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__9585 (
            .O(N__42543),
            .I(N__42540));
    LocalMux I__9584 (
            .O(N__42540),
            .I(N__42537));
    Span4Mux_h I__9583 (
            .O(N__42537),
            .I(N__42534));
    Odrv4 I__9582 (
            .O(N__42534),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__9581 (
            .O(N__42531),
            .I(N__42528));
    LocalMux I__9580 (
            .O(N__42528),
            .I(N__42525));
    Span4Mux_h I__9579 (
            .O(N__42525),
            .I(N__42522));
    Odrv4 I__9578 (
            .O(N__42522),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__9577 (
            .O(N__42519),
            .I(N__42516));
    LocalMux I__9576 (
            .O(N__42516),
            .I(N__42513));
    Span4Mux_h I__9575 (
            .O(N__42513),
            .I(N__42510));
    Odrv4 I__9574 (
            .O(N__42510),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__9573 (
            .O(N__42507),
            .I(N__42504));
    LocalMux I__9572 (
            .O(N__42504),
            .I(N__42501));
    Span4Mux_h I__9571 (
            .O(N__42501),
            .I(N__42498));
    Odrv4 I__9570 (
            .O(N__42498),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    CascadeMux I__9569 (
            .O(N__42495),
            .I(N__42492));
    InMux I__9568 (
            .O(N__42492),
            .I(N__42489));
    LocalMux I__9567 (
            .O(N__42489),
            .I(N__42484));
    InMux I__9566 (
            .O(N__42488),
            .I(N__42481));
    InMux I__9565 (
            .O(N__42487),
            .I(N__42478));
    Span4Mux_h I__9564 (
            .O(N__42484),
            .I(N__42473));
    LocalMux I__9563 (
            .O(N__42481),
            .I(N__42473));
    LocalMux I__9562 (
            .O(N__42478),
            .I(N__42469));
    Span4Mux_h I__9561 (
            .O(N__42473),
            .I(N__42466));
    InMux I__9560 (
            .O(N__42472),
            .I(N__42463));
    Odrv12 I__9559 (
            .O(N__42469),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__9558 (
            .O(N__42466),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__9557 (
            .O(N__42463),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__9556 (
            .O(N__42456),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__9555 (
            .O(N__42453),
            .I(N__42450));
    InMux I__9554 (
            .O(N__42450),
            .I(N__42446));
    InMux I__9553 (
            .O(N__42449),
            .I(N__42442));
    LocalMux I__9552 (
            .O(N__42446),
            .I(N__42439));
    InMux I__9551 (
            .O(N__42445),
            .I(N__42436));
    LocalMux I__9550 (
            .O(N__42442),
            .I(N__42431));
    Span4Mux_h I__9549 (
            .O(N__42439),
            .I(N__42431));
    LocalMux I__9548 (
            .O(N__42436),
            .I(N__42428));
    Span4Mux_h I__9547 (
            .O(N__42431),
            .I(N__42424));
    Span12Mux_h I__9546 (
            .O(N__42428),
            .I(N__42421));
    InMux I__9545 (
            .O(N__42427),
            .I(N__42418));
    Odrv4 I__9544 (
            .O(N__42424),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv12 I__9543 (
            .O(N__42421),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__9542 (
            .O(N__42418),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__9541 (
            .O(N__42411),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__9540 (
            .O(N__42408),
            .I(N__42404));
    InMux I__9539 (
            .O(N__42407),
            .I(N__42401));
    InMux I__9538 (
            .O(N__42404),
            .I(N__42396));
    LocalMux I__9537 (
            .O(N__42401),
            .I(N__42393));
    InMux I__9536 (
            .O(N__42400),
            .I(N__42390));
    InMux I__9535 (
            .O(N__42399),
            .I(N__42387));
    LocalMux I__9534 (
            .O(N__42396),
            .I(N__42382));
    Span4Mux_h I__9533 (
            .O(N__42393),
            .I(N__42382));
    LocalMux I__9532 (
            .O(N__42390),
            .I(N__42379));
    LocalMux I__9531 (
            .O(N__42387),
            .I(N__42374));
    Span4Mux_h I__9530 (
            .O(N__42382),
            .I(N__42374));
    Span4Mux_v I__9529 (
            .O(N__42379),
            .I(N__42371));
    Span4Mux_h I__9528 (
            .O(N__42374),
            .I(N__42368));
    Odrv4 I__9527 (
            .O(N__42371),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__9526 (
            .O(N__42368),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__9525 (
            .O(N__42363),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__9524 (
            .O(N__42360),
            .I(N__42356));
    CascadeMux I__9523 (
            .O(N__42359),
            .I(N__42353));
    InMux I__9522 (
            .O(N__42356),
            .I(N__42350));
    InMux I__9521 (
            .O(N__42353),
            .I(N__42347));
    LocalMux I__9520 (
            .O(N__42350),
            .I(N__42340));
    LocalMux I__9519 (
            .O(N__42347),
            .I(N__42340));
    InMux I__9518 (
            .O(N__42346),
            .I(N__42337));
    InMux I__9517 (
            .O(N__42345),
            .I(N__42334));
    Span4Mux_v I__9516 (
            .O(N__42340),
            .I(N__42327));
    LocalMux I__9515 (
            .O(N__42337),
            .I(N__42327));
    LocalMux I__9514 (
            .O(N__42334),
            .I(N__42327));
    Span4Mux_h I__9513 (
            .O(N__42327),
            .I(N__42324));
    Odrv4 I__9512 (
            .O(N__42324),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__9511 (
            .O(N__42321),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__9510 (
            .O(N__42318),
            .I(N__42315));
    InMux I__9509 (
            .O(N__42315),
            .I(N__42312));
    LocalMux I__9508 (
            .O(N__42312),
            .I(N__42309));
    Span4Mux_h I__9507 (
            .O(N__42309),
            .I(N__42306));
    Odrv4 I__9506 (
            .O(N__42306),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    InMux I__9505 (
            .O(N__42303),
            .I(N__42300));
    LocalMux I__9504 (
            .O(N__42300),
            .I(N__42297));
    Span4Mux_h I__9503 (
            .O(N__42297),
            .I(N__42293));
    InMux I__9502 (
            .O(N__42296),
            .I(N__42290));
    Odrv4 I__9501 (
            .O(N__42293),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    LocalMux I__9500 (
            .O(N__42290),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    InMux I__9499 (
            .O(N__42285),
            .I(N__42278));
    InMux I__9498 (
            .O(N__42284),
            .I(N__42278));
    InMux I__9497 (
            .O(N__42283),
            .I(N__42274));
    LocalMux I__9496 (
            .O(N__42278),
            .I(N__42271));
    InMux I__9495 (
            .O(N__42277),
            .I(N__42268));
    LocalMux I__9494 (
            .O(N__42274),
            .I(N__42263));
    Span4Mux_v I__9493 (
            .O(N__42271),
            .I(N__42263));
    LocalMux I__9492 (
            .O(N__42268),
            .I(N__42260));
    Odrv4 I__9491 (
            .O(N__42263),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    Odrv4 I__9490 (
            .O(N__42260),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    CascadeMux I__9489 (
            .O(N__42255),
            .I(elapsed_time_ns_1_RNI2COBB_0_15_cascade_));
    InMux I__9488 (
            .O(N__42252),
            .I(N__42249));
    LocalMux I__9487 (
            .O(N__42249),
            .I(N__42246));
    Odrv4 I__9486 (
            .O(N__42246),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__9485 (
            .O(N__42243),
            .I(N__42239));
    InMux I__9484 (
            .O(N__42242),
            .I(N__42236));
    LocalMux I__9483 (
            .O(N__42239),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    LocalMux I__9482 (
            .O(N__42236),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__9481 (
            .O(N__42231),
            .I(N__42226));
    InMux I__9480 (
            .O(N__42230),
            .I(N__42223));
    InMux I__9479 (
            .O(N__42229),
            .I(N__42220));
    LocalMux I__9478 (
            .O(N__42226),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__9477 (
            .O(N__42223),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__9476 (
            .O(N__42220),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    CascadeMux I__9475 (
            .O(N__42213),
            .I(N__42209));
    CascadeMux I__9474 (
            .O(N__42212),
            .I(N__42206));
    InMux I__9473 (
            .O(N__42209),
            .I(N__42203));
    InMux I__9472 (
            .O(N__42206),
            .I(N__42200));
    LocalMux I__9471 (
            .O(N__42203),
            .I(N__42195));
    LocalMux I__9470 (
            .O(N__42200),
            .I(N__42195));
    Odrv12 I__9469 (
            .O(N__42195),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__9468 (
            .O(N__42192),
            .I(N__42187));
    InMux I__9467 (
            .O(N__42191),
            .I(N__42184));
    InMux I__9466 (
            .O(N__42190),
            .I(N__42181));
    LocalMux I__9465 (
            .O(N__42187),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__9464 (
            .O(N__42184),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__9463 (
            .O(N__42181),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__9462 (
            .O(N__42174),
            .I(N__42171));
    LocalMux I__9461 (
            .O(N__42171),
            .I(N__42168));
    Span4Mux_h I__9460 (
            .O(N__42168),
            .I(N__42165));
    Odrv4 I__9459 (
            .O(N__42165),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__9458 (
            .O(N__42162),
            .I(N__42159));
    LocalMux I__9457 (
            .O(N__42159),
            .I(N__42156));
    Odrv12 I__9456 (
            .O(N__42156),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ));
    InMux I__9455 (
            .O(N__42153),
            .I(N__42150));
    LocalMux I__9454 (
            .O(N__42150),
            .I(N__42147));
    Odrv4 I__9453 (
            .O(N__42147),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__9452 (
            .O(N__42144),
            .I(N__42141));
    LocalMux I__9451 (
            .O(N__42141),
            .I(N__42138));
    Odrv4 I__9450 (
            .O(N__42138),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__9449 (
            .O(N__42135),
            .I(N__42132));
    LocalMux I__9448 (
            .O(N__42132),
            .I(N__42129));
    Span4Mux_v I__9447 (
            .O(N__42129),
            .I(N__42126));
    Odrv4 I__9446 (
            .O(N__42126),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    IoInMux I__9445 (
            .O(N__42123),
            .I(N__42089));
    InMux I__9444 (
            .O(N__42122),
            .I(N__42086));
    InMux I__9443 (
            .O(N__42121),
            .I(N__42079));
    InMux I__9442 (
            .O(N__42120),
            .I(N__42079));
    InMux I__9441 (
            .O(N__42119),
            .I(N__42079));
    InMux I__9440 (
            .O(N__42118),
            .I(N__42070));
    InMux I__9439 (
            .O(N__42117),
            .I(N__42070));
    InMux I__9438 (
            .O(N__42116),
            .I(N__42070));
    InMux I__9437 (
            .O(N__42115),
            .I(N__42070));
    InMux I__9436 (
            .O(N__42114),
            .I(N__42061));
    InMux I__9435 (
            .O(N__42113),
            .I(N__42061));
    InMux I__9434 (
            .O(N__42112),
            .I(N__42061));
    InMux I__9433 (
            .O(N__42111),
            .I(N__42061));
    InMux I__9432 (
            .O(N__42110),
            .I(N__42052));
    InMux I__9431 (
            .O(N__42109),
            .I(N__42052));
    InMux I__9430 (
            .O(N__42108),
            .I(N__42052));
    InMux I__9429 (
            .O(N__42107),
            .I(N__42052));
    InMux I__9428 (
            .O(N__42106),
            .I(N__42043));
    InMux I__9427 (
            .O(N__42105),
            .I(N__42043));
    InMux I__9426 (
            .O(N__42104),
            .I(N__42043));
    InMux I__9425 (
            .O(N__42103),
            .I(N__42043));
    InMux I__9424 (
            .O(N__42102),
            .I(N__42034));
    InMux I__9423 (
            .O(N__42101),
            .I(N__42034));
    InMux I__9422 (
            .O(N__42100),
            .I(N__42034));
    InMux I__9421 (
            .O(N__42099),
            .I(N__42034));
    InMux I__9420 (
            .O(N__42098),
            .I(N__42027));
    InMux I__9419 (
            .O(N__42097),
            .I(N__42027));
    InMux I__9418 (
            .O(N__42096),
            .I(N__42027));
    InMux I__9417 (
            .O(N__42095),
            .I(N__42018));
    InMux I__9416 (
            .O(N__42094),
            .I(N__42018));
    InMux I__9415 (
            .O(N__42093),
            .I(N__42018));
    InMux I__9414 (
            .O(N__42092),
            .I(N__42018));
    LocalMux I__9413 (
            .O(N__42089),
            .I(N__42015));
    LocalMux I__9412 (
            .O(N__42086),
            .I(N__42012));
    LocalMux I__9411 (
            .O(N__42079),
            .I(N__42007));
    LocalMux I__9410 (
            .O(N__42070),
            .I(N__42007));
    LocalMux I__9409 (
            .O(N__42061),
            .I(N__42002));
    LocalMux I__9408 (
            .O(N__42052),
            .I(N__42002));
    LocalMux I__9407 (
            .O(N__42043),
            .I(N__41997));
    LocalMux I__9406 (
            .O(N__42034),
            .I(N__41997));
    LocalMux I__9405 (
            .O(N__42027),
            .I(N__41992));
    LocalMux I__9404 (
            .O(N__42018),
            .I(N__41992));
    IoSpan4Mux I__9403 (
            .O(N__42015),
            .I(N__41989));
    Span4Mux_h I__9402 (
            .O(N__42012),
            .I(N__41984));
    Span4Mux_h I__9401 (
            .O(N__42007),
            .I(N__41984));
    Span4Mux_h I__9400 (
            .O(N__42002),
            .I(N__41981));
    Span4Mux_h I__9399 (
            .O(N__41997),
            .I(N__41978));
    Span12Mux_s10_h I__9398 (
            .O(N__41992),
            .I(N__41975));
    Span4Mux_s1_v I__9397 (
            .O(N__41989),
            .I(N__41970));
    Span4Mux_v I__9396 (
            .O(N__41984),
            .I(N__41970));
    Span4Mux_v I__9395 (
            .O(N__41981),
            .I(N__41967));
    Odrv4 I__9394 (
            .O(N__41978),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv12 I__9393 (
            .O(N__41975),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__9392 (
            .O(N__41970),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__9391 (
            .O(N__41967),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__9390 (
            .O(N__41958),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__9389 (
            .O(N__41955),
            .I(N__41952));
    LocalMux I__9388 (
            .O(N__41952),
            .I(N__41948));
    CascadeMux I__9387 (
            .O(N__41951),
            .I(N__41945));
    Span4Mux_h I__9386 (
            .O(N__41948),
            .I(N__41941));
    InMux I__9385 (
            .O(N__41945),
            .I(N__41937));
    InMux I__9384 (
            .O(N__41944),
            .I(N__41934));
    Sp12to4 I__9383 (
            .O(N__41941),
            .I(N__41931));
    InMux I__9382 (
            .O(N__41940),
            .I(N__41928));
    LocalMux I__9381 (
            .O(N__41937),
            .I(N__41924));
    LocalMux I__9380 (
            .O(N__41934),
            .I(N__41921));
    Span12Mux_v I__9379 (
            .O(N__41931),
            .I(N__41918));
    LocalMux I__9378 (
            .O(N__41928),
            .I(N__41915));
    InMux I__9377 (
            .O(N__41927),
            .I(N__41912));
    Span4Mux_v I__9376 (
            .O(N__41924),
            .I(N__41909));
    Span12Mux_v I__9375 (
            .O(N__41921),
            .I(N__41904));
    Span12Mux_v I__9374 (
            .O(N__41918),
            .I(N__41904));
    Span4Mux_h I__9373 (
            .O(N__41915),
            .I(N__41901));
    LocalMux I__9372 (
            .O(N__41912),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__9371 (
            .O(N__41909),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv12 I__9370 (
            .O(N__41904),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__9369 (
            .O(N__41901),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    IoInMux I__9368 (
            .O(N__41892),
            .I(N__41889));
    LocalMux I__9367 (
            .O(N__41889),
            .I(N__41886));
    Span12Mux_s8_v I__9366 (
            .O(N__41886),
            .I(N__41883));
    Span12Mux_v I__9365 (
            .O(N__41883),
            .I(N__41879));
    InMux I__9364 (
            .O(N__41882),
            .I(N__41876));
    Odrv12 I__9363 (
            .O(N__41879),
            .I(T23_c));
    LocalMux I__9362 (
            .O(N__41876),
            .I(T23_c));
    InMux I__9361 (
            .O(N__41871),
            .I(N__41868));
    LocalMux I__9360 (
            .O(N__41868),
            .I(N__41864));
    InMux I__9359 (
            .O(N__41867),
            .I(N__41861));
    Span4Mux_v I__9358 (
            .O(N__41864),
            .I(N__41858));
    LocalMux I__9357 (
            .O(N__41861),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    Odrv4 I__9356 (
            .O(N__41858),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    CascadeMux I__9355 (
            .O(N__41853),
            .I(N__41850));
    InMux I__9354 (
            .O(N__41850),
            .I(N__41847));
    LocalMux I__9353 (
            .O(N__41847),
            .I(N__41844));
    Span4Mux_v I__9352 (
            .O(N__41844),
            .I(N__41841));
    Odrv4 I__9351 (
            .O(N__41841),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df30 ));
    InMux I__9350 (
            .O(N__41838),
            .I(N__41835));
    LocalMux I__9349 (
            .O(N__41835),
            .I(N__41829));
    InMux I__9348 (
            .O(N__41834),
            .I(N__41824));
    InMux I__9347 (
            .O(N__41833),
            .I(N__41824));
    InMux I__9346 (
            .O(N__41832),
            .I(N__41821));
    Span4Mux_v I__9345 (
            .O(N__41829),
            .I(N__41818));
    LocalMux I__9344 (
            .O(N__41824),
            .I(N__41815));
    LocalMux I__9343 (
            .O(N__41821),
            .I(N__41812));
    Odrv4 I__9342 (
            .O(N__41818),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__9341 (
            .O(N__41815),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__9340 (
            .O(N__41812),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__9339 (
            .O(N__41805),
            .I(N__41802));
    LocalMux I__9338 (
            .O(N__41802),
            .I(N__41799));
    Span4Mux_v I__9337 (
            .O(N__41799),
            .I(N__41795));
    InMux I__9336 (
            .O(N__41798),
            .I(N__41792));
    Odrv4 I__9335 (
            .O(N__41795),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    LocalMux I__9334 (
            .O(N__41792),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    InMux I__9333 (
            .O(N__41787),
            .I(N__41778));
    InMux I__9332 (
            .O(N__41786),
            .I(N__41778));
    InMux I__9331 (
            .O(N__41785),
            .I(N__41778));
    LocalMux I__9330 (
            .O(N__41778),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    InMux I__9329 (
            .O(N__41775),
            .I(N__41769));
    InMux I__9328 (
            .O(N__41774),
            .I(N__41762));
    InMux I__9327 (
            .O(N__41773),
            .I(N__41762));
    InMux I__9326 (
            .O(N__41772),
            .I(N__41762));
    LocalMux I__9325 (
            .O(N__41769),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__9324 (
            .O(N__41762),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    CascadeMux I__9323 (
            .O(N__41757),
            .I(N__41752));
    CascadeMux I__9322 (
            .O(N__41756),
            .I(N__41749));
    InMux I__9321 (
            .O(N__41755),
            .I(N__41745));
    InMux I__9320 (
            .O(N__41752),
            .I(N__41738));
    InMux I__9319 (
            .O(N__41749),
            .I(N__41738));
    InMux I__9318 (
            .O(N__41748),
            .I(N__41738));
    LocalMux I__9317 (
            .O(N__41745),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__9316 (
            .O(N__41738),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    CascadeMux I__9315 (
            .O(N__41733),
            .I(N__41730));
    InMux I__9314 (
            .O(N__41730),
            .I(N__41727));
    LocalMux I__9313 (
            .O(N__41727),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    CascadeMux I__9312 (
            .O(N__41724),
            .I(N__41720));
    InMux I__9311 (
            .O(N__41723),
            .I(N__41712));
    InMux I__9310 (
            .O(N__41720),
            .I(N__41712));
    InMux I__9309 (
            .O(N__41719),
            .I(N__41712));
    LocalMux I__9308 (
            .O(N__41712),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    InMux I__9307 (
            .O(N__41709),
            .I(N__41704));
    InMux I__9306 (
            .O(N__41708),
            .I(N__41699));
    InMux I__9305 (
            .O(N__41707),
            .I(N__41699));
    LocalMux I__9304 (
            .O(N__41704),
            .I(N__41693));
    LocalMux I__9303 (
            .O(N__41699),
            .I(N__41693));
    InMux I__9302 (
            .O(N__41698),
            .I(N__41690));
    Span4Mux_h I__9301 (
            .O(N__41693),
            .I(N__41685));
    LocalMux I__9300 (
            .O(N__41690),
            .I(N__41685));
    Odrv4 I__9299 (
            .O(N__41685),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__9298 (
            .O(N__41682),
            .I(N__41679));
    LocalMux I__9297 (
            .O(N__41679),
            .I(N__41675));
    InMux I__9296 (
            .O(N__41678),
            .I(N__41672));
    Odrv4 I__9295 (
            .O(N__41675),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    LocalMux I__9294 (
            .O(N__41672),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    InMux I__9293 (
            .O(N__41667),
            .I(N__41664));
    LocalMux I__9292 (
            .O(N__41664),
            .I(N__41661));
    Odrv4 I__9291 (
            .O(N__41661),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    InMux I__9290 (
            .O(N__41658),
            .I(N__41651));
    InMux I__9289 (
            .O(N__41657),
            .I(N__41651));
    InMux I__9288 (
            .O(N__41656),
            .I(N__41648));
    LocalMux I__9287 (
            .O(N__41651),
            .I(N__41645));
    LocalMux I__9286 (
            .O(N__41648),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__9285 (
            .O(N__41645),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__9284 (
            .O(N__41640),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    CascadeMux I__9283 (
            .O(N__41637),
            .I(N__41634));
    InMux I__9282 (
            .O(N__41634),
            .I(N__41627));
    InMux I__9281 (
            .O(N__41633),
            .I(N__41627));
    InMux I__9280 (
            .O(N__41632),
            .I(N__41624));
    LocalMux I__9279 (
            .O(N__41627),
            .I(N__41621));
    LocalMux I__9278 (
            .O(N__41624),
            .I(N__41616));
    Span4Mux_v I__9277 (
            .O(N__41621),
            .I(N__41616));
    Odrv4 I__9276 (
            .O(N__41616),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__9275 (
            .O(N__41613),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__9274 (
            .O(N__41610),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__9273 (
            .O(N__41607),
            .I(bfn_17_10_0_));
    InMux I__9272 (
            .O(N__41604),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__9271 (
            .O(N__41601),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__9270 (
            .O(N__41598),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__9269 (
            .O(N__41595),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__9268 (
            .O(N__41592),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__9267 (
            .O(N__41589),
            .I(N__41585));
    InMux I__9266 (
            .O(N__41588),
            .I(N__41582));
    LocalMux I__9265 (
            .O(N__41585),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__9264 (
            .O(N__41582),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__9263 (
            .O(N__41577),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__9262 (
            .O(N__41574),
            .I(N__41570));
    InMux I__9261 (
            .O(N__41573),
            .I(N__41567));
    LocalMux I__9260 (
            .O(N__41570),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__9259 (
            .O(N__41567),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__9258 (
            .O(N__41562),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__9257 (
            .O(N__41559),
            .I(N__41555));
    InMux I__9256 (
            .O(N__41558),
            .I(N__41552));
    LocalMux I__9255 (
            .O(N__41555),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__9254 (
            .O(N__41552),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__9253 (
            .O(N__41547),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__9252 (
            .O(N__41544),
            .I(N__41537));
    InMux I__9251 (
            .O(N__41543),
            .I(N__41537));
    InMux I__9250 (
            .O(N__41542),
            .I(N__41534));
    LocalMux I__9249 (
            .O(N__41537),
            .I(N__41531));
    LocalMux I__9248 (
            .O(N__41534),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__9247 (
            .O(N__41531),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__9246 (
            .O(N__41526),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    CascadeMux I__9245 (
            .O(N__41523),
            .I(N__41519));
    InMux I__9244 (
            .O(N__41522),
            .I(N__41514));
    InMux I__9243 (
            .O(N__41519),
            .I(N__41514));
    LocalMux I__9242 (
            .O(N__41514),
            .I(N__41510));
    InMux I__9241 (
            .O(N__41513),
            .I(N__41507));
    Span4Mux_v I__9240 (
            .O(N__41510),
            .I(N__41504));
    LocalMux I__9239 (
            .O(N__41507),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__9238 (
            .O(N__41504),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__9237 (
            .O(N__41499),
            .I(bfn_17_9_0_));
    InMux I__9236 (
            .O(N__41496),
            .I(N__41489));
    InMux I__9235 (
            .O(N__41495),
            .I(N__41489));
    InMux I__9234 (
            .O(N__41494),
            .I(N__41486));
    LocalMux I__9233 (
            .O(N__41489),
            .I(N__41483));
    LocalMux I__9232 (
            .O(N__41486),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__9231 (
            .O(N__41483),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__9230 (
            .O(N__41478),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    CascadeMux I__9229 (
            .O(N__41475),
            .I(N__41472));
    InMux I__9228 (
            .O(N__41472),
            .I(N__41465));
    InMux I__9227 (
            .O(N__41471),
            .I(N__41465));
    InMux I__9226 (
            .O(N__41470),
            .I(N__41462));
    LocalMux I__9225 (
            .O(N__41465),
            .I(N__41459));
    LocalMux I__9224 (
            .O(N__41462),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__9223 (
            .O(N__41459),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__9222 (
            .O(N__41454),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__9221 (
            .O(N__41451),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__9220 (
            .O(N__41448),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__9219 (
            .O(N__41445),
            .I(N__41441));
    InMux I__9218 (
            .O(N__41444),
            .I(N__41438));
    LocalMux I__9217 (
            .O(N__41441),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__9216 (
            .O(N__41438),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__9215 (
            .O(N__41433),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__9214 (
            .O(N__41430),
            .I(N__41427));
    LocalMux I__9213 (
            .O(N__41427),
            .I(N__41423));
    InMux I__9212 (
            .O(N__41426),
            .I(N__41420));
    Span4Mux_v I__9211 (
            .O(N__41423),
            .I(N__41417));
    LocalMux I__9210 (
            .O(N__41420),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__9209 (
            .O(N__41417),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__9208 (
            .O(N__41412),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__9207 (
            .O(N__41409),
            .I(N__41405));
    InMux I__9206 (
            .O(N__41408),
            .I(N__41402));
    LocalMux I__9205 (
            .O(N__41405),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__9204 (
            .O(N__41402),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__9203 (
            .O(N__41397),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__9202 (
            .O(N__41394),
            .I(N__41390));
    InMux I__9201 (
            .O(N__41393),
            .I(N__41387));
    LocalMux I__9200 (
            .O(N__41390),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__9199 (
            .O(N__41387),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__9198 (
            .O(N__41382),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__9197 (
            .O(N__41379),
            .I(N__41375));
    InMux I__9196 (
            .O(N__41378),
            .I(N__41372));
    LocalMux I__9195 (
            .O(N__41375),
            .I(N__41369));
    LocalMux I__9194 (
            .O(N__41372),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__9193 (
            .O(N__41369),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__9192 (
            .O(N__41364),
            .I(bfn_17_8_0_));
    InMux I__9191 (
            .O(N__41361),
            .I(N__41357));
    InMux I__9190 (
            .O(N__41360),
            .I(N__41354));
    LocalMux I__9189 (
            .O(N__41357),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__9188 (
            .O(N__41354),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__9187 (
            .O(N__41349),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__9186 (
            .O(N__41346),
            .I(N__41342));
    InMux I__9185 (
            .O(N__41345),
            .I(N__41339));
    LocalMux I__9184 (
            .O(N__41342),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__9183 (
            .O(N__41339),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__9182 (
            .O(N__41334),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__9181 (
            .O(N__41331),
            .I(N__41327));
    InMux I__9180 (
            .O(N__41330),
            .I(N__41324));
    LocalMux I__9179 (
            .O(N__41327),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__9178 (
            .O(N__41324),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__9177 (
            .O(N__41319),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__9176 (
            .O(N__41316),
            .I(N__41313));
    LocalMux I__9175 (
            .O(N__41313),
            .I(N__41310));
    Odrv4 I__9174 (
            .O(N__41310),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__9173 (
            .O(N__41307),
            .I(N__41303));
    InMux I__9172 (
            .O(N__41306),
            .I(N__41298));
    LocalMux I__9171 (
            .O(N__41303),
            .I(N__41295));
    InMux I__9170 (
            .O(N__41302),
            .I(N__41290));
    InMux I__9169 (
            .O(N__41301),
            .I(N__41290));
    LocalMux I__9168 (
            .O(N__41298),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__9167 (
            .O(N__41295),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__9166 (
            .O(N__41290),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__9165 (
            .O(N__41283),
            .I(N__41274));
    InMux I__9164 (
            .O(N__41282),
            .I(N__41274));
    InMux I__9163 (
            .O(N__41281),
            .I(N__41271));
    InMux I__9162 (
            .O(N__41280),
            .I(N__41266));
    InMux I__9161 (
            .O(N__41279),
            .I(N__41266));
    LocalMux I__9160 (
            .O(N__41274),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__9159 (
            .O(N__41271),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__9158 (
            .O(N__41266),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__9157 (
            .O(N__41259),
            .I(N__41255));
    InMux I__9156 (
            .O(N__41258),
            .I(N__41252));
    LocalMux I__9155 (
            .O(N__41255),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__9154 (
            .O(N__41252),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    InMux I__9153 (
            .O(N__41247),
            .I(N__41244));
    LocalMux I__9152 (
            .O(N__41244),
            .I(N__41239));
    InMux I__9151 (
            .O(N__41243),
            .I(N__41236));
    InMux I__9150 (
            .O(N__41242),
            .I(N__41232));
    Span4Mux_v I__9149 (
            .O(N__41239),
            .I(N__41229));
    LocalMux I__9148 (
            .O(N__41236),
            .I(N__41226));
    InMux I__9147 (
            .O(N__41235),
            .I(N__41223));
    LocalMux I__9146 (
            .O(N__41232),
            .I(N__41220));
    Sp12to4 I__9145 (
            .O(N__41229),
            .I(N__41217));
    Span4Mux_h I__9144 (
            .O(N__41226),
            .I(N__41212));
    LocalMux I__9143 (
            .O(N__41223),
            .I(N__41212));
    Span4Mux_h I__9142 (
            .O(N__41220),
            .I(N__41209));
    Span12Mux_h I__9141 (
            .O(N__41217),
            .I(N__41206));
    Span4Mux_h I__9140 (
            .O(N__41212),
            .I(N__41203));
    Odrv4 I__9139 (
            .O(N__41209),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv12 I__9138 (
            .O(N__41206),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__9137 (
            .O(N__41203),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__9136 (
            .O(N__41196),
            .I(N__41193));
    LocalMux I__9135 (
            .O(N__41193),
            .I(N__41156));
    InMux I__9134 (
            .O(N__41192),
            .I(N__41147));
    InMux I__9133 (
            .O(N__41191),
            .I(N__41147));
    InMux I__9132 (
            .O(N__41190),
            .I(N__41147));
    InMux I__9131 (
            .O(N__41189),
            .I(N__41147));
    InMux I__9130 (
            .O(N__41188),
            .I(N__41144));
    CascadeMux I__9129 (
            .O(N__41187),
            .I(N__41139));
    InMux I__9128 (
            .O(N__41186),
            .I(N__41129));
    CascadeMux I__9127 (
            .O(N__41185),
            .I(N__41116));
    InMux I__9126 (
            .O(N__41184),
            .I(N__41112));
    InMux I__9125 (
            .O(N__41183),
            .I(N__41106));
    InMux I__9124 (
            .O(N__41182),
            .I(N__41099));
    InMux I__9123 (
            .O(N__41181),
            .I(N__41099));
    InMux I__9122 (
            .O(N__41180),
            .I(N__41087));
    InMux I__9121 (
            .O(N__41179),
            .I(N__41087));
    InMux I__9120 (
            .O(N__41178),
            .I(N__41078));
    InMux I__9119 (
            .O(N__41177),
            .I(N__41078));
    InMux I__9118 (
            .O(N__41176),
            .I(N__41078));
    InMux I__9117 (
            .O(N__41175),
            .I(N__41078));
    InMux I__9116 (
            .O(N__41174),
            .I(N__41069));
    InMux I__9115 (
            .O(N__41173),
            .I(N__41069));
    InMux I__9114 (
            .O(N__41172),
            .I(N__41069));
    InMux I__9113 (
            .O(N__41171),
            .I(N__41069));
    InMux I__9112 (
            .O(N__41170),
            .I(N__41066));
    InMux I__9111 (
            .O(N__41169),
            .I(N__41063));
    InMux I__9110 (
            .O(N__41168),
            .I(N__41060));
    InMux I__9109 (
            .O(N__41167),
            .I(N__41057));
    InMux I__9108 (
            .O(N__41166),
            .I(N__41050));
    InMux I__9107 (
            .O(N__41165),
            .I(N__41050));
    InMux I__9106 (
            .O(N__41164),
            .I(N__41050));
    InMux I__9105 (
            .O(N__41163),
            .I(N__41045));
    InMux I__9104 (
            .O(N__41162),
            .I(N__41045));
    InMux I__9103 (
            .O(N__41161),
            .I(N__41038));
    InMux I__9102 (
            .O(N__41160),
            .I(N__41038));
    InMux I__9101 (
            .O(N__41159),
            .I(N__41038));
    Span4Mux_h I__9100 (
            .O(N__41156),
            .I(N__41031));
    LocalMux I__9099 (
            .O(N__41147),
            .I(N__41031));
    LocalMux I__9098 (
            .O(N__41144),
            .I(N__41031));
    InMux I__9097 (
            .O(N__41143),
            .I(N__41024));
    InMux I__9096 (
            .O(N__41142),
            .I(N__41024));
    InMux I__9095 (
            .O(N__41139),
            .I(N__41024));
    InMux I__9094 (
            .O(N__41138),
            .I(N__41021));
    InMux I__9093 (
            .O(N__41137),
            .I(N__41018));
    InMux I__9092 (
            .O(N__41136),
            .I(N__41011));
    InMux I__9091 (
            .O(N__41135),
            .I(N__41011));
    InMux I__9090 (
            .O(N__41134),
            .I(N__41011));
    InMux I__9089 (
            .O(N__41133),
            .I(N__41006));
    InMux I__9088 (
            .O(N__41132),
            .I(N__41006));
    LocalMux I__9087 (
            .O(N__41129),
            .I(N__41003));
    InMux I__9086 (
            .O(N__41128),
            .I(N__40973));
    InMux I__9085 (
            .O(N__41127),
            .I(N__40973));
    InMux I__9084 (
            .O(N__41126),
            .I(N__40973));
    InMux I__9083 (
            .O(N__41125),
            .I(N__40973));
    InMux I__9082 (
            .O(N__41124),
            .I(N__40973));
    InMux I__9081 (
            .O(N__41123),
            .I(N__40973));
    InMux I__9080 (
            .O(N__41122),
            .I(N__40973));
    InMux I__9079 (
            .O(N__41121),
            .I(N__40973));
    InMux I__9078 (
            .O(N__41120),
            .I(N__40964));
    InMux I__9077 (
            .O(N__41119),
            .I(N__40964));
    InMux I__9076 (
            .O(N__41116),
            .I(N__40964));
    InMux I__9075 (
            .O(N__41115),
            .I(N__40964));
    LocalMux I__9074 (
            .O(N__41112),
            .I(N__40961));
    CascadeMux I__9073 (
            .O(N__41111),
            .I(N__40958));
    InMux I__9072 (
            .O(N__41110),
            .I(N__40941));
    InMux I__9071 (
            .O(N__41109),
            .I(N__40941));
    LocalMux I__9070 (
            .O(N__41106),
            .I(N__40938));
    InMux I__9069 (
            .O(N__41105),
            .I(N__40933));
    InMux I__9068 (
            .O(N__41104),
            .I(N__40933));
    LocalMux I__9067 (
            .O(N__41099),
            .I(N__40930));
    InMux I__9066 (
            .O(N__41098),
            .I(N__40919));
    InMux I__9065 (
            .O(N__41097),
            .I(N__40919));
    InMux I__9064 (
            .O(N__41096),
            .I(N__40919));
    InMux I__9063 (
            .O(N__41095),
            .I(N__40919));
    InMux I__9062 (
            .O(N__41094),
            .I(N__40919));
    InMux I__9061 (
            .O(N__41093),
            .I(N__40914));
    InMux I__9060 (
            .O(N__41092),
            .I(N__40914));
    LocalMux I__9059 (
            .O(N__41087),
            .I(N__40905));
    LocalMux I__9058 (
            .O(N__41078),
            .I(N__40905));
    LocalMux I__9057 (
            .O(N__41069),
            .I(N__40905));
    LocalMux I__9056 (
            .O(N__41066),
            .I(N__40905));
    LocalMux I__9055 (
            .O(N__41063),
            .I(N__40902));
    LocalMux I__9054 (
            .O(N__41060),
            .I(N__40899));
    LocalMux I__9053 (
            .O(N__41057),
            .I(N__40886));
    LocalMux I__9052 (
            .O(N__41050),
            .I(N__40886));
    LocalMux I__9051 (
            .O(N__41045),
            .I(N__40886));
    LocalMux I__9050 (
            .O(N__41038),
            .I(N__40886));
    Span4Mux_v I__9049 (
            .O(N__41031),
            .I(N__40886));
    LocalMux I__9048 (
            .O(N__41024),
            .I(N__40886));
    LocalMux I__9047 (
            .O(N__41021),
            .I(N__40881));
    LocalMux I__9046 (
            .O(N__41018),
            .I(N__40881));
    LocalMux I__9045 (
            .O(N__41011),
            .I(N__40876));
    LocalMux I__9044 (
            .O(N__41006),
            .I(N__40876));
    Span4Mux_v I__9043 (
            .O(N__41003),
            .I(N__40873));
    InMux I__9042 (
            .O(N__41002),
            .I(N__40870));
    InMux I__9041 (
            .O(N__41001),
            .I(N__40857));
    InMux I__9040 (
            .O(N__41000),
            .I(N__40857));
    InMux I__9039 (
            .O(N__40999),
            .I(N__40857));
    InMux I__9038 (
            .O(N__40998),
            .I(N__40857));
    InMux I__9037 (
            .O(N__40997),
            .I(N__40857));
    InMux I__9036 (
            .O(N__40996),
            .I(N__40857));
    InMux I__9035 (
            .O(N__40995),
            .I(N__40844));
    InMux I__9034 (
            .O(N__40994),
            .I(N__40844));
    InMux I__9033 (
            .O(N__40993),
            .I(N__40844));
    InMux I__9032 (
            .O(N__40992),
            .I(N__40844));
    InMux I__9031 (
            .O(N__40991),
            .I(N__40844));
    InMux I__9030 (
            .O(N__40990),
            .I(N__40844));
    LocalMux I__9029 (
            .O(N__40973),
            .I(N__40837));
    LocalMux I__9028 (
            .O(N__40964),
            .I(N__40837));
    Span4Mux_h I__9027 (
            .O(N__40961),
            .I(N__40837));
    InMux I__9026 (
            .O(N__40958),
            .I(N__40828));
    InMux I__9025 (
            .O(N__40957),
            .I(N__40828));
    InMux I__9024 (
            .O(N__40956),
            .I(N__40828));
    InMux I__9023 (
            .O(N__40955),
            .I(N__40828));
    InMux I__9022 (
            .O(N__40954),
            .I(N__40821));
    InMux I__9021 (
            .O(N__40953),
            .I(N__40821));
    InMux I__9020 (
            .O(N__40952),
            .I(N__40821));
    InMux I__9019 (
            .O(N__40951),
            .I(N__40814));
    InMux I__9018 (
            .O(N__40950),
            .I(N__40814));
    InMux I__9017 (
            .O(N__40949),
            .I(N__40814));
    InMux I__9016 (
            .O(N__40948),
            .I(N__40807));
    InMux I__9015 (
            .O(N__40947),
            .I(N__40807));
    InMux I__9014 (
            .O(N__40946),
            .I(N__40807));
    LocalMux I__9013 (
            .O(N__40941),
            .I(N__40798));
    Span4Mux_v I__9012 (
            .O(N__40938),
            .I(N__40798));
    LocalMux I__9011 (
            .O(N__40933),
            .I(N__40798));
    Span4Mux_h I__9010 (
            .O(N__40930),
            .I(N__40798));
    LocalMux I__9009 (
            .O(N__40919),
            .I(N__40789));
    LocalMux I__9008 (
            .O(N__40914),
            .I(N__40789));
    Sp12to4 I__9007 (
            .O(N__40905),
            .I(N__40789));
    Span12Mux_s10_h I__9006 (
            .O(N__40902),
            .I(N__40789));
    Span4Mux_v I__9005 (
            .O(N__40899),
            .I(N__40778));
    Span4Mux_v I__9004 (
            .O(N__40886),
            .I(N__40778));
    Span4Mux_v I__9003 (
            .O(N__40881),
            .I(N__40778));
    Span4Mux_h I__9002 (
            .O(N__40876),
            .I(N__40778));
    Span4Mux_h I__9001 (
            .O(N__40873),
            .I(N__40778));
    LocalMux I__9000 (
            .O(N__40870),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8999 (
            .O(N__40857),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8998 (
            .O(N__40844),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__8997 (
            .O(N__40837),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8996 (
            .O(N__40828),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8995 (
            .O(N__40821),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8994 (
            .O(N__40814),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8993 (
            .O(N__40807),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__8992 (
            .O(N__40798),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__8991 (
            .O(N__40789),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__8990 (
            .O(N__40778),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__8989 (
            .O(N__40755),
            .I(N__40752));
    LocalMux I__8988 (
            .O(N__40752),
            .I(N__40748));
    InMux I__8987 (
            .O(N__40751),
            .I(N__40745));
    Span4Mux_h I__8986 (
            .O(N__40748),
            .I(N__40742));
    LocalMux I__8985 (
            .O(N__40745),
            .I(N__40739));
    Span4Mux_h I__8984 (
            .O(N__40742),
            .I(N__40735));
    Span4Mux_h I__8983 (
            .O(N__40739),
            .I(N__40732));
    InMux I__8982 (
            .O(N__40738),
            .I(N__40729));
    Span4Mux_v I__8981 (
            .O(N__40735),
            .I(N__40726));
    Span4Mux_h I__8980 (
            .O(N__40732),
            .I(N__40723));
    LocalMux I__8979 (
            .O(N__40729),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    Odrv4 I__8978 (
            .O(N__40726),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    Odrv4 I__8977 (
            .O(N__40723),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    CascadeMux I__8976 (
            .O(N__40716),
            .I(N__40712));
    InMux I__8975 (
            .O(N__40715),
            .I(N__40708));
    InMux I__8974 (
            .O(N__40712),
            .I(N__40705));
    InMux I__8973 (
            .O(N__40711),
            .I(N__40702));
    LocalMux I__8972 (
            .O(N__40708),
            .I(N__40699));
    LocalMux I__8971 (
            .O(N__40705),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__8970 (
            .O(N__40702),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__8969 (
            .O(N__40699),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__8968 (
            .O(N__40692),
            .I(N__40689));
    InMux I__8967 (
            .O(N__40689),
            .I(N__40686));
    LocalMux I__8966 (
            .O(N__40686),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    InMux I__8965 (
            .O(N__40683),
            .I(N__40679));
    InMux I__8964 (
            .O(N__40682),
            .I(N__40676));
    LocalMux I__8963 (
            .O(N__40679),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__8962 (
            .O(N__40676),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__8961 (
            .O(N__40671),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__8960 (
            .O(N__40668),
            .I(N__40665));
    LocalMux I__8959 (
            .O(N__40665),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ));
    CascadeMux I__8958 (
            .O(N__40662),
            .I(N__40659));
    InMux I__8957 (
            .O(N__40659),
            .I(N__40655));
    InMux I__8956 (
            .O(N__40658),
            .I(N__40652));
    LocalMux I__8955 (
            .O(N__40655),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__8954 (
            .O(N__40652),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__8953 (
            .O(N__40647),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__8952 (
            .O(N__40644),
            .I(N__40640));
    InMux I__8951 (
            .O(N__40643),
            .I(N__40637));
    LocalMux I__8950 (
            .O(N__40640),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__8949 (
            .O(N__40637),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__8948 (
            .O(N__40632),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__8947 (
            .O(N__40629),
            .I(N__40622));
    CascadeMux I__8946 (
            .O(N__40628),
            .I(N__40618));
    CascadeMux I__8945 (
            .O(N__40627),
            .I(N__40591));
    CascadeMux I__8944 (
            .O(N__40626),
            .I(N__40588));
    InMux I__8943 (
            .O(N__40625),
            .I(N__40567));
    LocalMux I__8942 (
            .O(N__40622),
            .I(N__40561));
    InMux I__8941 (
            .O(N__40621),
            .I(N__40544));
    InMux I__8940 (
            .O(N__40618),
            .I(N__40544));
    InMux I__8939 (
            .O(N__40617),
            .I(N__40544));
    InMux I__8938 (
            .O(N__40616),
            .I(N__40544));
    InMux I__8937 (
            .O(N__40615),
            .I(N__40544));
    InMux I__8936 (
            .O(N__40614),
            .I(N__40544));
    InMux I__8935 (
            .O(N__40613),
            .I(N__40544));
    InMux I__8934 (
            .O(N__40612),
            .I(N__40544));
    InMux I__8933 (
            .O(N__40611),
            .I(N__40531));
    InMux I__8932 (
            .O(N__40610),
            .I(N__40531));
    InMux I__8931 (
            .O(N__40609),
            .I(N__40531));
    InMux I__8930 (
            .O(N__40608),
            .I(N__40531));
    InMux I__8929 (
            .O(N__40607),
            .I(N__40531));
    InMux I__8928 (
            .O(N__40606),
            .I(N__40531));
    InMux I__8927 (
            .O(N__40605),
            .I(N__40528));
    InMux I__8926 (
            .O(N__40604),
            .I(N__40519));
    InMux I__8925 (
            .O(N__40603),
            .I(N__40519));
    InMux I__8924 (
            .O(N__40602),
            .I(N__40519));
    InMux I__8923 (
            .O(N__40601),
            .I(N__40519));
    InMux I__8922 (
            .O(N__40600),
            .I(N__40512));
    InMux I__8921 (
            .O(N__40599),
            .I(N__40512));
    InMux I__8920 (
            .O(N__40598),
            .I(N__40512));
    InMux I__8919 (
            .O(N__40597),
            .I(N__40507));
    InMux I__8918 (
            .O(N__40596),
            .I(N__40507));
    InMux I__8917 (
            .O(N__40595),
            .I(N__40502));
    InMux I__8916 (
            .O(N__40594),
            .I(N__40502));
    InMux I__8915 (
            .O(N__40591),
            .I(N__40487));
    InMux I__8914 (
            .O(N__40588),
            .I(N__40487));
    InMux I__8913 (
            .O(N__40587),
            .I(N__40487));
    InMux I__8912 (
            .O(N__40586),
            .I(N__40487));
    InMux I__8911 (
            .O(N__40585),
            .I(N__40487));
    InMux I__8910 (
            .O(N__40584),
            .I(N__40487));
    InMux I__8909 (
            .O(N__40583),
            .I(N__40487));
    InMux I__8908 (
            .O(N__40582),
            .I(N__40479));
    InMux I__8907 (
            .O(N__40581),
            .I(N__40476));
    InMux I__8906 (
            .O(N__40580),
            .I(N__40473));
    InMux I__8905 (
            .O(N__40579),
            .I(N__40466));
    InMux I__8904 (
            .O(N__40578),
            .I(N__40466));
    InMux I__8903 (
            .O(N__40577),
            .I(N__40466));
    InMux I__8902 (
            .O(N__40576),
            .I(N__40453));
    InMux I__8901 (
            .O(N__40575),
            .I(N__40453));
    InMux I__8900 (
            .O(N__40574),
            .I(N__40453));
    InMux I__8899 (
            .O(N__40573),
            .I(N__40453));
    InMux I__8898 (
            .O(N__40572),
            .I(N__40453));
    InMux I__8897 (
            .O(N__40571),
            .I(N__40453));
    InMux I__8896 (
            .O(N__40570),
            .I(N__40438));
    LocalMux I__8895 (
            .O(N__40567),
            .I(N__40435));
    InMux I__8894 (
            .O(N__40566),
            .I(N__40428));
    InMux I__8893 (
            .O(N__40565),
            .I(N__40428));
    InMux I__8892 (
            .O(N__40564),
            .I(N__40428));
    Span4Mux_h I__8891 (
            .O(N__40561),
            .I(N__40423));
    LocalMux I__8890 (
            .O(N__40544),
            .I(N__40423));
    LocalMux I__8889 (
            .O(N__40531),
            .I(N__40420));
    LocalMux I__8888 (
            .O(N__40528),
            .I(N__40417));
    LocalMux I__8887 (
            .O(N__40519),
            .I(N__40412));
    LocalMux I__8886 (
            .O(N__40512),
            .I(N__40412));
    LocalMux I__8885 (
            .O(N__40507),
            .I(N__40407));
    LocalMux I__8884 (
            .O(N__40502),
            .I(N__40407));
    LocalMux I__8883 (
            .O(N__40487),
            .I(N__40404));
    InMux I__8882 (
            .O(N__40486),
            .I(N__40393));
    InMux I__8881 (
            .O(N__40485),
            .I(N__40393));
    InMux I__8880 (
            .O(N__40484),
            .I(N__40393));
    InMux I__8879 (
            .O(N__40483),
            .I(N__40393));
    InMux I__8878 (
            .O(N__40482),
            .I(N__40393));
    LocalMux I__8877 (
            .O(N__40479),
            .I(N__40388));
    LocalMux I__8876 (
            .O(N__40476),
            .I(N__40388));
    LocalMux I__8875 (
            .O(N__40473),
            .I(N__40381));
    LocalMux I__8874 (
            .O(N__40466),
            .I(N__40381));
    LocalMux I__8873 (
            .O(N__40453),
            .I(N__40381));
    InMux I__8872 (
            .O(N__40452),
            .I(N__40364));
    InMux I__8871 (
            .O(N__40451),
            .I(N__40364));
    InMux I__8870 (
            .O(N__40450),
            .I(N__40364));
    InMux I__8869 (
            .O(N__40449),
            .I(N__40364));
    InMux I__8868 (
            .O(N__40448),
            .I(N__40364));
    InMux I__8867 (
            .O(N__40447),
            .I(N__40364));
    InMux I__8866 (
            .O(N__40446),
            .I(N__40364));
    InMux I__8865 (
            .O(N__40445),
            .I(N__40364));
    InMux I__8864 (
            .O(N__40444),
            .I(N__40358));
    InMux I__8863 (
            .O(N__40443),
            .I(N__40351));
    InMux I__8862 (
            .O(N__40442),
            .I(N__40351));
    InMux I__8861 (
            .O(N__40441),
            .I(N__40351));
    LocalMux I__8860 (
            .O(N__40438),
            .I(N__40344));
    Span4Mux_v I__8859 (
            .O(N__40435),
            .I(N__40344));
    LocalMux I__8858 (
            .O(N__40428),
            .I(N__40344));
    Span4Mux_v I__8857 (
            .O(N__40423),
            .I(N__40339));
    Span4Mux_h I__8856 (
            .O(N__40420),
            .I(N__40339));
    Span4Mux_v I__8855 (
            .O(N__40417),
            .I(N__40336));
    Span4Mux_v I__8854 (
            .O(N__40412),
            .I(N__40333));
    Span4Mux_h I__8853 (
            .O(N__40407),
            .I(N__40326));
    Span4Mux_h I__8852 (
            .O(N__40404),
            .I(N__40326));
    LocalMux I__8851 (
            .O(N__40393),
            .I(N__40326));
    Span4Mux_h I__8850 (
            .O(N__40388),
            .I(N__40319));
    Span4Mux_v I__8849 (
            .O(N__40381),
            .I(N__40319));
    LocalMux I__8848 (
            .O(N__40364),
            .I(N__40319));
    InMux I__8847 (
            .O(N__40363),
            .I(N__40312));
    InMux I__8846 (
            .O(N__40362),
            .I(N__40312));
    InMux I__8845 (
            .O(N__40361),
            .I(N__40312));
    LocalMux I__8844 (
            .O(N__40358),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__8843 (
            .O(N__40351),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__8842 (
            .O(N__40344),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__8841 (
            .O(N__40339),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__8840 (
            .O(N__40336),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__8839 (
            .O(N__40333),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__8838 (
            .O(N__40326),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__8837 (
            .O(N__40319),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__8836 (
            .O(N__40312),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__8835 (
            .O(N__40293),
            .I(N__40288));
    InMux I__8834 (
            .O(N__40292),
            .I(N__40285));
    InMux I__8833 (
            .O(N__40291),
            .I(N__40282));
    LocalMux I__8832 (
            .O(N__40288),
            .I(N__40279));
    LocalMux I__8831 (
            .O(N__40285),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__8830 (
            .O(N__40282),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv12 I__8829 (
            .O(N__40279),
            .I(\current_shift_inst.un4_control_input1_27 ));
    CascadeMux I__8828 (
            .O(N__40272),
            .I(N__40257));
    CascadeMux I__8827 (
            .O(N__40271),
            .I(N__40253));
    CascadeMux I__8826 (
            .O(N__40270),
            .I(N__40250));
    CascadeMux I__8825 (
            .O(N__40269),
            .I(N__40247));
    CascadeMux I__8824 (
            .O(N__40268),
            .I(N__40242));
    CascadeMux I__8823 (
            .O(N__40267),
            .I(N__40239));
    CascadeMux I__8822 (
            .O(N__40266),
            .I(N__40225));
    InMux I__8821 (
            .O(N__40265),
            .I(N__40218));
    InMux I__8820 (
            .O(N__40264),
            .I(N__40218));
    InMux I__8819 (
            .O(N__40263),
            .I(N__40218));
    InMux I__8818 (
            .O(N__40262),
            .I(N__40209));
    InMux I__8817 (
            .O(N__40261),
            .I(N__40209));
    InMux I__8816 (
            .O(N__40260),
            .I(N__40209));
    InMux I__8815 (
            .O(N__40257),
            .I(N__40209));
    CascadeMux I__8814 (
            .O(N__40256),
            .I(N__40205));
    InMux I__8813 (
            .O(N__40253),
            .I(N__40192));
    InMux I__8812 (
            .O(N__40250),
            .I(N__40187));
    InMux I__8811 (
            .O(N__40247),
            .I(N__40187));
    InMux I__8810 (
            .O(N__40246),
            .I(N__40182));
    InMux I__8809 (
            .O(N__40245),
            .I(N__40182));
    InMux I__8808 (
            .O(N__40242),
            .I(N__40179));
    InMux I__8807 (
            .O(N__40239),
            .I(N__40176));
    CascadeMux I__8806 (
            .O(N__40238),
            .I(N__40171));
    CascadeMux I__8805 (
            .O(N__40237),
            .I(N__40167));
    CascadeMux I__8804 (
            .O(N__40236),
            .I(N__40164));
    CascadeMux I__8803 (
            .O(N__40235),
            .I(N__40160));
    CascadeMux I__8802 (
            .O(N__40234),
            .I(N__40157));
    CascadeMux I__8801 (
            .O(N__40233),
            .I(N__40154));
    CascadeMux I__8800 (
            .O(N__40232),
            .I(N__40151));
    CascadeMux I__8799 (
            .O(N__40231),
            .I(N__40147));
    CascadeMux I__8798 (
            .O(N__40230),
            .I(N__40130));
    CascadeMux I__8797 (
            .O(N__40229),
            .I(N__40122));
    InMux I__8796 (
            .O(N__40228),
            .I(N__40115));
    InMux I__8795 (
            .O(N__40225),
            .I(N__40115));
    LocalMux I__8794 (
            .O(N__40218),
            .I(N__40106));
    LocalMux I__8793 (
            .O(N__40209),
            .I(N__40106));
    InMux I__8792 (
            .O(N__40208),
            .I(N__40101));
    InMux I__8791 (
            .O(N__40205),
            .I(N__40101));
    InMux I__8790 (
            .O(N__40204),
            .I(N__40086));
    InMux I__8789 (
            .O(N__40203),
            .I(N__40086));
    InMux I__8788 (
            .O(N__40202),
            .I(N__40086));
    InMux I__8787 (
            .O(N__40201),
            .I(N__40086));
    InMux I__8786 (
            .O(N__40200),
            .I(N__40086));
    InMux I__8785 (
            .O(N__40199),
            .I(N__40086));
    InMux I__8784 (
            .O(N__40198),
            .I(N__40086));
    InMux I__8783 (
            .O(N__40197),
            .I(N__40079));
    InMux I__8782 (
            .O(N__40196),
            .I(N__40079));
    InMux I__8781 (
            .O(N__40195),
            .I(N__40079));
    LocalMux I__8780 (
            .O(N__40192),
            .I(N__40076));
    LocalMux I__8779 (
            .O(N__40187),
            .I(N__40073));
    LocalMux I__8778 (
            .O(N__40182),
            .I(N__40066));
    LocalMux I__8777 (
            .O(N__40179),
            .I(N__40066));
    LocalMux I__8776 (
            .O(N__40176),
            .I(N__40066));
    InMux I__8775 (
            .O(N__40175),
            .I(N__40061));
    InMux I__8774 (
            .O(N__40174),
            .I(N__40061));
    InMux I__8773 (
            .O(N__40171),
            .I(N__40052));
    InMux I__8772 (
            .O(N__40170),
            .I(N__40052));
    InMux I__8771 (
            .O(N__40167),
            .I(N__40052));
    InMux I__8770 (
            .O(N__40164),
            .I(N__40052));
    InMux I__8769 (
            .O(N__40163),
            .I(N__40043));
    InMux I__8768 (
            .O(N__40160),
            .I(N__40043));
    InMux I__8767 (
            .O(N__40157),
            .I(N__40043));
    InMux I__8766 (
            .O(N__40154),
            .I(N__40043));
    InMux I__8765 (
            .O(N__40151),
            .I(N__40040));
    InMux I__8764 (
            .O(N__40150),
            .I(N__40035));
    InMux I__8763 (
            .O(N__40147),
            .I(N__40035));
    CascadeMux I__8762 (
            .O(N__40146),
            .I(N__40030));
    CascadeMux I__8761 (
            .O(N__40145),
            .I(N__40026));
    CascadeMux I__8760 (
            .O(N__40144),
            .I(N__40022));
    CascadeMux I__8759 (
            .O(N__40143),
            .I(N__40017));
    CascadeMux I__8758 (
            .O(N__40142),
            .I(N__40013));
    CascadeMux I__8757 (
            .O(N__40141),
            .I(N__40009));
    CascadeMux I__8756 (
            .O(N__40140),
            .I(N__40004));
    CascadeMux I__8755 (
            .O(N__40139),
            .I(N__40000));
    CascadeMux I__8754 (
            .O(N__40138),
            .I(N__39996));
    CascadeMux I__8753 (
            .O(N__40137),
            .I(N__39992));
    CascadeMux I__8752 (
            .O(N__40136),
            .I(N__39989));
    CascadeMux I__8751 (
            .O(N__40135),
            .I(N__39985));
    CascadeMux I__8750 (
            .O(N__40134),
            .I(N__39981));
    CascadeMux I__8749 (
            .O(N__40133),
            .I(N__39977));
    InMux I__8748 (
            .O(N__40130),
            .I(N__39962));
    CascadeMux I__8747 (
            .O(N__40129),
            .I(N__39959));
    InMux I__8746 (
            .O(N__40128),
            .I(N__39939));
    InMux I__8745 (
            .O(N__40127),
            .I(N__39939));
    InMux I__8744 (
            .O(N__40126),
            .I(N__39939));
    InMux I__8743 (
            .O(N__40125),
            .I(N__39939));
    InMux I__8742 (
            .O(N__40122),
            .I(N__39939));
    InMux I__8741 (
            .O(N__40121),
            .I(N__39939));
    InMux I__8740 (
            .O(N__40120),
            .I(N__39939));
    LocalMux I__8739 (
            .O(N__40115),
            .I(N__39936));
    InMux I__8738 (
            .O(N__40114),
            .I(N__39927));
    InMux I__8737 (
            .O(N__40113),
            .I(N__39927));
    InMux I__8736 (
            .O(N__40112),
            .I(N__39927));
    InMux I__8735 (
            .O(N__40111),
            .I(N__39927));
    Span4Mux_v I__8734 (
            .O(N__40106),
            .I(N__39918));
    LocalMux I__8733 (
            .O(N__40101),
            .I(N__39918));
    LocalMux I__8732 (
            .O(N__40086),
            .I(N__39918));
    LocalMux I__8731 (
            .O(N__40079),
            .I(N__39918));
    Span4Mux_v I__8730 (
            .O(N__40076),
            .I(N__39901));
    Span4Mux_h I__8729 (
            .O(N__40073),
            .I(N__39901));
    Span4Mux_v I__8728 (
            .O(N__40066),
            .I(N__39901));
    LocalMux I__8727 (
            .O(N__40061),
            .I(N__39901));
    LocalMux I__8726 (
            .O(N__40052),
            .I(N__39901));
    LocalMux I__8725 (
            .O(N__40043),
            .I(N__39901));
    LocalMux I__8724 (
            .O(N__40040),
            .I(N__39901));
    LocalMux I__8723 (
            .O(N__40035),
            .I(N__39901));
    InMux I__8722 (
            .O(N__40034),
            .I(N__39884));
    InMux I__8721 (
            .O(N__40033),
            .I(N__39884));
    InMux I__8720 (
            .O(N__40030),
            .I(N__39884));
    InMux I__8719 (
            .O(N__40029),
            .I(N__39884));
    InMux I__8718 (
            .O(N__40026),
            .I(N__39884));
    InMux I__8717 (
            .O(N__40025),
            .I(N__39884));
    InMux I__8716 (
            .O(N__40022),
            .I(N__39884));
    InMux I__8715 (
            .O(N__40021),
            .I(N__39884));
    InMux I__8714 (
            .O(N__40020),
            .I(N__39869));
    InMux I__8713 (
            .O(N__40017),
            .I(N__39869));
    InMux I__8712 (
            .O(N__40016),
            .I(N__39869));
    InMux I__8711 (
            .O(N__40013),
            .I(N__39869));
    InMux I__8710 (
            .O(N__40012),
            .I(N__39869));
    InMux I__8709 (
            .O(N__40009),
            .I(N__39869));
    InMux I__8708 (
            .O(N__40008),
            .I(N__39869));
    InMux I__8707 (
            .O(N__40007),
            .I(N__39852));
    InMux I__8706 (
            .O(N__40004),
            .I(N__39852));
    InMux I__8705 (
            .O(N__40003),
            .I(N__39852));
    InMux I__8704 (
            .O(N__40000),
            .I(N__39852));
    InMux I__8703 (
            .O(N__39999),
            .I(N__39852));
    InMux I__8702 (
            .O(N__39996),
            .I(N__39852));
    InMux I__8701 (
            .O(N__39995),
            .I(N__39852));
    InMux I__8700 (
            .O(N__39992),
            .I(N__39852));
    InMux I__8699 (
            .O(N__39989),
            .I(N__39835));
    InMux I__8698 (
            .O(N__39988),
            .I(N__39835));
    InMux I__8697 (
            .O(N__39985),
            .I(N__39835));
    InMux I__8696 (
            .O(N__39984),
            .I(N__39835));
    InMux I__8695 (
            .O(N__39981),
            .I(N__39835));
    InMux I__8694 (
            .O(N__39980),
            .I(N__39835));
    InMux I__8693 (
            .O(N__39977),
            .I(N__39835));
    InMux I__8692 (
            .O(N__39976),
            .I(N__39835));
    CascadeMux I__8691 (
            .O(N__39975),
            .I(N__39832));
    CascadeMux I__8690 (
            .O(N__39974),
            .I(N__39828));
    CascadeMux I__8689 (
            .O(N__39973),
            .I(N__39824));
    CascadeMux I__8688 (
            .O(N__39972),
            .I(N__39820));
    CascadeMux I__8687 (
            .O(N__39971),
            .I(N__39816));
    CascadeMux I__8686 (
            .O(N__39970),
            .I(N__39812));
    CascadeMux I__8685 (
            .O(N__39969),
            .I(N__39808));
    CascadeMux I__8684 (
            .O(N__39968),
            .I(N__39804));
    CascadeMux I__8683 (
            .O(N__39967),
            .I(N__39796));
    CascadeMux I__8682 (
            .O(N__39966),
            .I(N__39792));
    CascadeMux I__8681 (
            .O(N__39965),
            .I(N__39788));
    LocalMux I__8680 (
            .O(N__39962),
            .I(N__39782));
    InMux I__8679 (
            .O(N__39959),
            .I(N__39779));
    InMux I__8678 (
            .O(N__39958),
            .I(N__39768));
    InMux I__8677 (
            .O(N__39957),
            .I(N__39768));
    InMux I__8676 (
            .O(N__39956),
            .I(N__39768));
    InMux I__8675 (
            .O(N__39955),
            .I(N__39768));
    InMux I__8674 (
            .O(N__39954),
            .I(N__39768));
    LocalMux I__8673 (
            .O(N__39939),
            .I(N__39765));
    Span4Mux_h I__8672 (
            .O(N__39936),
            .I(N__39758));
    LocalMux I__8671 (
            .O(N__39927),
            .I(N__39758));
    Span4Mux_v I__8670 (
            .O(N__39918),
            .I(N__39758));
    Span4Mux_h I__8669 (
            .O(N__39901),
            .I(N__39747));
    LocalMux I__8668 (
            .O(N__39884),
            .I(N__39747));
    LocalMux I__8667 (
            .O(N__39869),
            .I(N__39747));
    LocalMux I__8666 (
            .O(N__39852),
            .I(N__39747));
    LocalMux I__8665 (
            .O(N__39835),
            .I(N__39747));
    InMux I__8664 (
            .O(N__39832),
            .I(N__39730));
    InMux I__8663 (
            .O(N__39831),
            .I(N__39730));
    InMux I__8662 (
            .O(N__39828),
            .I(N__39730));
    InMux I__8661 (
            .O(N__39827),
            .I(N__39730));
    InMux I__8660 (
            .O(N__39824),
            .I(N__39730));
    InMux I__8659 (
            .O(N__39823),
            .I(N__39730));
    InMux I__8658 (
            .O(N__39820),
            .I(N__39730));
    InMux I__8657 (
            .O(N__39819),
            .I(N__39730));
    InMux I__8656 (
            .O(N__39816),
            .I(N__39713));
    InMux I__8655 (
            .O(N__39815),
            .I(N__39713));
    InMux I__8654 (
            .O(N__39812),
            .I(N__39713));
    InMux I__8653 (
            .O(N__39811),
            .I(N__39713));
    InMux I__8652 (
            .O(N__39808),
            .I(N__39713));
    InMux I__8651 (
            .O(N__39807),
            .I(N__39713));
    InMux I__8650 (
            .O(N__39804),
            .I(N__39713));
    InMux I__8649 (
            .O(N__39803),
            .I(N__39713));
    InMux I__8648 (
            .O(N__39802),
            .I(N__39706));
    InMux I__8647 (
            .O(N__39801),
            .I(N__39706));
    InMux I__8646 (
            .O(N__39800),
            .I(N__39706));
    InMux I__8645 (
            .O(N__39799),
            .I(N__39693));
    InMux I__8644 (
            .O(N__39796),
            .I(N__39693));
    InMux I__8643 (
            .O(N__39795),
            .I(N__39693));
    InMux I__8642 (
            .O(N__39792),
            .I(N__39693));
    InMux I__8641 (
            .O(N__39791),
            .I(N__39693));
    InMux I__8640 (
            .O(N__39788),
            .I(N__39693));
    InMux I__8639 (
            .O(N__39787),
            .I(N__39686));
    InMux I__8638 (
            .O(N__39786),
            .I(N__39686));
    InMux I__8637 (
            .O(N__39785),
            .I(N__39686));
    Odrv4 I__8636 (
            .O(N__39782),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__8635 (
            .O(N__39779),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__8634 (
            .O(N__39768),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__8633 (
            .O(N__39765),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__8632 (
            .O(N__39758),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__8631 (
            .O(N__39747),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__8630 (
            .O(N__39730),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__8629 (
            .O(N__39713),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__8628 (
            .O(N__39706),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__8627 (
            .O(N__39693),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__8626 (
            .O(N__39686),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__8625 (
            .O(N__39663),
            .I(N__39660));
    InMux I__8624 (
            .O(N__39660),
            .I(N__39657));
    LocalMux I__8623 (
            .O(N__39657),
            .I(N__39654));
    Span4Mux_v I__8622 (
            .O(N__39654),
            .I(N__39651));
    Span4Mux_h I__8621 (
            .O(N__39651),
            .I(N__39648));
    Odrv4 I__8620 (
            .O(N__39648),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__8619 (
            .O(N__39645),
            .I(N__39642));
    LocalMux I__8618 (
            .O(N__39642),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__8617 (
            .O(N__39639),
            .I(N__39636));
    LocalMux I__8616 (
            .O(N__39636),
            .I(N__39633));
    Odrv4 I__8615 (
            .O(N__39633),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__8614 (
            .O(N__39630),
            .I(N__39627));
    LocalMux I__8613 (
            .O(N__39627),
            .I(N__39624));
    Odrv4 I__8612 (
            .O(N__39624),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__8611 (
            .O(N__39621),
            .I(N__39618));
    LocalMux I__8610 (
            .O(N__39618),
            .I(N__39615));
    Odrv4 I__8609 (
            .O(N__39615),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__8608 (
            .O(N__39612),
            .I(N__39609));
    LocalMux I__8607 (
            .O(N__39609),
            .I(N__39606));
    Odrv4 I__8606 (
            .O(N__39606),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__8605 (
            .O(N__39603),
            .I(N__39600));
    LocalMux I__8604 (
            .O(N__39600),
            .I(N__39596));
    InMux I__8603 (
            .O(N__39599),
            .I(N__39593));
    Span4Mux_h I__8602 (
            .O(N__39596),
            .I(N__39590));
    LocalMux I__8601 (
            .O(N__39593),
            .I(N__39587));
    Span4Mux_v I__8600 (
            .O(N__39590),
            .I(N__39584));
    Span4Mux_v I__8599 (
            .O(N__39587),
            .I(N__39580));
    Span4Mux_v I__8598 (
            .O(N__39584),
            .I(N__39577));
    CascadeMux I__8597 (
            .O(N__39583),
            .I(N__39572));
    Span4Mux_v I__8596 (
            .O(N__39580),
            .I(N__39569));
    Span4Mux_v I__8595 (
            .O(N__39577),
            .I(N__39566));
    InMux I__8594 (
            .O(N__39576),
            .I(N__39563));
    InMux I__8593 (
            .O(N__39575),
            .I(N__39560));
    InMux I__8592 (
            .O(N__39572),
            .I(N__39557));
    Span4Mux_v I__8591 (
            .O(N__39569),
            .I(N__39554));
    Span4Mux_v I__8590 (
            .O(N__39566),
            .I(N__39551));
    LocalMux I__8589 (
            .O(N__39563),
            .I(N__39548));
    LocalMux I__8588 (
            .O(N__39560),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__8587 (
            .O(N__39557),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__8586 (
            .O(N__39554),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__8585 (
            .O(N__39551),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__8584 (
            .O(N__39548),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    IoInMux I__8583 (
            .O(N__39537),
            .I(N__39534));
    LocalMux I__8582 (
            .O(N__39534),
            .I(N__39531));
    Span12Mux_s1_v I__8581 (
            .O(N__39531),
            .I(N__39528));
    Span12Mux_v I__8580 (
            .O(N__39528),
            .I(N__39524));
    InMux I__8579 (
            .O(N__39527),
            .I(N__39521));
    Odrv12 I__8578 (
            .O(N__39524),
            .I(T01_c));
    LocalMux I__8577 (
            .O(N__39521),
            .I(T01_c));
    InMux I__8576 (
            .O(N__39516),
            .I(N__39513));
    LocalMux I__8575 (
            .O(N__39513),
            .I(N__39510));
    Odrv4 I__8574 (
            .O(N__39510),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__8573 (
            .O(N__39507),
            .I(N__39504));
    LocalMux I__8572 (
            .O(N__39504),
            .I(N__39501));
    Odrv4 I__8571 (
            .O(N__39501),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__8570 (
            .O(N__39498),
            .I(N__39494));
    InMux I__8569 (
            .O(N__39497),
            .I(N__39491));
    LocalMux I__8568 (
            .O(N__39494),
            .I(N__39487));
    LocalMux I__8567 (
            .O(N__39491),
            .I(N__39484));
    InMux I__8566 (
            .O(N__39490),
            .I(N__39481));
    Span4Mux_h I__8565 (
            .O(N__39487),
            .I(N__39477));
    Span4Mux_h I__8564 (
            .O(N__39484),
            .I(N__39472));
    LocalMux I__8563 (
            .O(N__39481),
            .I(N__39472));
    InMux I__8562 (
            .O(N__39480),
            .I(N__39469));
    Odrv4 I__8561 (
            .O(N__39477),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    Odrv4 I__8560 (
            .O(N__39472),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__8559 (
            .O(N__39469),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__8558 (
            .O(N__39462),
            .I(N__39459));
    LocalMux I__8557 (
            .O(N__39459),
            .I(N__39456));
    Odrv4 I__8556 (
            .O(N__39456),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    InMux I__8555 (
            .O(N__39453),
            .I(N__39449));
    CascadeMux I__8554 (
            .O(N__39452),
            .I(N__39446));
    LocalMux I__8553 (
            .O(N__39449),
            .I(N__39441));
    InMux I__8552 (
            .O(N__39446),
            .I(N__39438));
    InMux I__8551 (
            .O(N__39445),
            .I(N__39432));
    InMux I__8550 (
            .O(N__39444),
            .I(N__39432));
    Span4Mux_v I__8549 (
            .O(N__39441),
            .I(N__39429));
    LocalMux I__8548 (
            .O(N__39438),
            .I(N__39426));
    InMux I__8547 (
            .O(N__39437),
            .I(N__39423));
    LocalMux I__8546 (
            .O(N__39432),
            .I(N__39420));
    Odrv4 I__8545 (
            .O(N__39429),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv12 I__8544 (
            .O(N__39426),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__8543 (
            .O(N__39423),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__8542 (
            .O(N__39420),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__8541 (
            .O(N__39411),
            .I(N__39408));
    LocalMux I__8540 (
            .O(N__39408),
            .I(N__39403));
    InMux I__8539 (
            .O(N__39407),
            .I(N__39400));
    InMux I__8538 (
            .O(N__39406),
            .I(N__39397));
    Span4Mux_v I__8537 (
            .O(N__39403),
            .I(N__39394));
    LocalMux I__8536 (
            .O(N__39400),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    LocalMux I__8535 (
            .O(N__39397),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv4 I__8534 (
            .O(N__39394),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__8533 (
            .O(N__39387),
            .I(N__39384));
    InMux I__8532 (
            .O(N__39384),
            .I(N__39381));
    LocalMux I__8531 (
            .O(N__39381),
            .I(N__39378));
    Span4Mux_v I__8530 (
            .O(N__39378),
            .I(N__39375));
    Span4Mux_h I__8529 (
            .O(N__39375),
            .I(N__39372));
    Odrv4 I__8528 (
            .O(N__39372),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__8527 (
            .O(N__39369),
            .I(N__39366));
    LocalMux I__8526 (
            .O(N__39366),
            .I(N__39361));
    InMux I__8525 (
            .O(N__39365),
            .I(N__39358));
    InMux I__8524 (
            .O(N__39364),
            .I(N__39355));
    Span4Mux_v I__8523 (
            .O(N__39361),
            .I(N__39350));
    LocalMux I__8522 (
            .O(N__39358),
            .I(N__39350));
    LocalMux I__8521 (
            .O(N__39355),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__8520 (
            .O(N__39350),
            .I(\current_shift_inst.un4_control_input1_23 ));
    CascadeMux I__8519 (
            .O(N__39345),
            .I(N__39342));
    InMux I__8518 (
            .O(N__39342),
            .I(N__39339));
    LocalMux I__8517 (
            .O(N__39339),
            .I(N__39336));
    Sp12to4 I__8516 (
            .O(N__39336),
            .I(N__39333));
    Span12Mux_v I__8515 (
            .O(N__39333),
            .I(N__39330));
    Odrv12 I__8514 (
            .O(N__39330),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__8513 (
            .O(N__39327),
            .I(N__39324));
    LocalMux I__8512 (
            .O(N__39324),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__8511 (
            .O(N__39321),
            .I(N__39318));
    LocalMux I__8510 (
            .O(N__39318),
            .I(N__39315));
    Odrv4 I__8509 (
            .O(N__39315),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__8508 (
            .O(N__39312),
            .I(N__39309));
    LocalMux I__8507 (
            .O(N__39309),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__8506 (
            .O(N__39306),
            .I(N__39303));
    LocalMux I__8505 (
            .O(N__39303),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__8504 (
            .O(N__39300),
            .I(N__39297));
    LocalMux I__8503 (
            .O(N__39297),
            .I(N__39294));
    Odrv4 I__8502 (
            .O(N__39294),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__8501 (
            .O(N__39291),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__8500 (
            .O(N__39288),
            .I(bfn_16_14_0_));
    InMux I__8499 (
            .O(N__39285),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__8498 (
            .O(N__39282),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__8497 (
            .O(N__39279),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__8496 (
            .O(N__39276),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    CascadeMux I__8495 (
            .O(N__39273),
            .I(N__39268));
    CascadeMux I__8494 (
            .O(N__39272),
            .I(N__39265));
    InMux I__8493 (
            .O(N__39271),
            .I(N__39258));
    InMux I__8492 (
            .O(N__39268),
            .I(N__39258));
    InMux I__8491 (
            .O(N__39265),
            .I(N__39258));
    LocalMux I__8490 (
            .O(N__39258),
            .I(N__39254));
    InMux I__8489 (
            .O(N__39257),
            .I(N__39251));
    Span4Mux_h I__8488 (
            .O(N__39254),
            .I(N__39248));
    LocalMux I__8487 (
            .O(N__39251),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__8486 (
            .O(N__39248),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__8485 (
            .O(N__39243),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__8484 (
            .O(N__39240),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    CascadeMux I__8483 (
            .O(N__39237),
            .I(N__39234));
    InMux I__8482 (
            .O(N__39234),
            .I(N__39225));
    InMux I__8481 (
            .O(N__39233),
            .I(N__39225));
    InMux I__8480 (
            .O(N__39232),
            .I(N__39225));
    LocalMux I__8479 (
            .O(N__39225),
            .I(N__39221));
    InMux I__8478 (
            .O(N__39224),
            .I(N__39218));
    Span4Mux_v I__8477 (
            .O(N__39221),
            .I(N__39215));
    LocalMux I__8476 (
            .O(N__39218),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__8475 (
            .O(N__39215),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__8474 (
            .O(N__39210),
            .I(N__39207));
    LocalMux I__8473 (
            .O(N__39207),
            .I(N__39203));
    InMux I__8472 (
            .O(N__39206),
            .I(N__39200));
    Span4Mux_h I__8471 (
            .O(N__39203),
            .I(N__39197));
    LocalMux I__8470 (
            .O(N__39200),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__8469 (
            .O(N__39197),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__8468 (
            .O(N__39192),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    CascadeMux I__8467 (
            .O(N__39189),
            .I(N__39186));
    InMux I__8466 (
            .O(N__39186),
            .I(N__39179));
    InMux I__8465 (
            .O(N__39185),
            .I(N__39179));
    InMux I__8464 (
            .O(N__39184),
            .I(N__39176));
    LocalMux I__8463 (
            .O(N__39179),
            .I(N__39173));
    LocalMux I__8462 (
            .O(N__39176),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__8461 (
            .O(N__39173),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__8460 (
            .O(N__39168),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__8459 (
            .O(N__39165),
            .I(N__39158));
    InMux I__8458 (
            .O(N__39164),
            .I(N__39158));
    InMux I__8457 (
            .O(N__39163),
            .I(N__39155));
    LocalMux I__8456 (
            .O(N__39158),
            .I(N__39152));
    LocalMux I__8455 (
            .O(N__39155),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__8454 (
            .O(N__39152),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__8453 (
            .O(N__39147),
            .I(bfn_16_13_0_));
    InMux I__8452 (
            .O(N__39144),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__8451 (
            .O(N__39141),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    CascadeMux I__8450 (
            .O(N__39138),
            .I(N__39134));
    InMux I__8449 (
            .O(N__39137),
            .I(N__39128));
    InMux I__8448 (
            .O(N__39134),
            .I(N__39128));
    InMux I__8447 (
            .O(N__39133),
            .I(N__39125));
    LocalMux I__8446 (
            .O(N__39128),
            .I(N__39122));
    LocalMux I__8445 (
            .O(N__39125),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__8444 (
            .O(N__39122),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__8443 (
            .O(N__39117),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__8442 (
            .O(N__39114),
            .I(N__39107));
    InMux I__8441 (
            .O(N__39113),
            .I(N__39107));
    InMux I__8440 (
            .O(N__39112),
            .I(N__39104));
    LocalMux I__8439 (
            .O(N__39107),
            .I(N__39101));
    LocalMux I__8438 (
            .O(N__39104),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__8437 (
            .O(N__39101),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__8436 (
            .O(N__39096),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__8435 (
            .O(N__39093),
            .I(N__39090));
    InMux I__8434 (
            .O(N__39090),
            .I(N__39084));
    InMux I__8433 (
            .O(N__39089),
            .I(N__39084));
    LocalMux I__8432 (
            .O(N__39084),
            .I(N__39080));
    InMux I__8431 (
            .O(N__39083),
            .I(N__39077));
    Span4Mux_h I__8430 (
            .O(N__39080),
            .I(N__39074));
    LocalMux I__8429 (
            .O(N__39077),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__8428 (
            .O(N__39074),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__8427 (
            .O(N__39069),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__8426 (
            .O(N__39066),
            .I(N__39060));
    InMux I__8425 (
            .O(N__39065),
            .I(N__39060));
    LocalMux I__8424 (
            .O(N__39060),
            .I(N__39056));
    InMux I__8423 (
            .O(N__39059),
            .I(N__39053));
    Span4Mux_h I__8422 (
            .O(N__39056),
            .I(N__39050));
    LocalMux I__8421 (
            .O(N__39053),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__8420 (
            .O(N__39050),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__8419 (
            .O(N__39045),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__8418 (
            .O(N__39042),
            .I(N__39038));
    InMux I__8417 (
            .O(N__39041),
            .I(N__39035));
    LocalMux I__8416 (
            .O(N__39038),
            .I(N__39032));
    LocalMux I__8415 (
            .O(N__39035),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__8414 (
            .O(N__39032),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__8413 (
            .O(N__39027),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__8412 (
            .O(N__39024),
            .I(N__39020));
    InMux I__8411 (
            .O(N__39023),
            .I(N__39017));
    LocalMux I__8410 (
            .O(N__39020),
            .I(N__39014));
    LocalMux I__8409 (
            .O(N__39017),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__8408 (
            .O(N__39014),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__8407 (
            .O(N__39009),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__8406 (
            .O(N__39006),
            .I(N__39002));
    InMux I__8405 (
            .O(N__39005),
            .I(N__38999));
    LocalMux I__8404 (
            .O(N__39002),
            .I(N__38996));
    LocalMux I__8403 (
            .O(N__38999),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__8402 (
            .O(N__38996),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__8401 (
            .O(N__38991),
            .I(bfn_16_12_0_));
    InMux I__8400 (
            .O(N__38988),
            .I(N__38984));
    InMux I__8399 (
            .O(N__38987),
            .I(N__38981));
    LocalMux I__8398 (
            .O(N__38984),
            .I(N__38978));
    LocalMux I__8397 (
            .O(N__38981),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__8396 (
            .O(N__38978),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__8395 (
            .O(N__38973),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__8394 (
            .O(N__38970),
            .I(N__38966));
    InMux I__8393 (
            .O(N__38969),
            .I(N__38963));
    LocalMux I__8392 (
            .O(N__38966),
            .I(N__38960));
    LocalMux I__8391 (
            .O(N__38963),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__8390 (
            .O(N__38960),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__8389 (
            .O(N__38955),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__8388 (
            .O(N__38952),
            .I(N__38948));
    InMux I__8387 (
            .O(N__38951),
            .I(N__38945));
    LocalMux I__8386 (
            .O(N__38948),
            .I(N__38942));
    LocalMux I__8385 (
            .O(N__38945),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__8384 (
            .O(N__38942),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__8383 (
            .O(N__38937),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__8382 (
            .O(N__38934),
            .I(N__38930));
    InMux I__8381 (
            .O(N__38933),
            .I(N__38927));
    LocalMux I__8380 (
            .O(N__38930),
            .I(N__38924));
    LocalMux I__8379 (
            .O(N__38927),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__8378 (
            .O(N__38924),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__8377 (
            .O(N__38919),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__8376 (
            .O(N__38916),
            .I(N__38912));
    InMux I__8375 (
            .O(N__38915),
            .I(N__38909));
    LocalMux I__8374 (
            .O(N__38912),
            .I(N__38906));
    LocalMux I__8373 (
            .O(N__38909),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv12 I__8372 (
            .O(N__38906),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__8371 (
            .O(N__38901),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__8370 (
            .O(N__38898),
            .I(N__38895));
    LocalMux I__8369 (
            .O(N__38895),
            .I(N__38892));
    Odrv12 I__8368 (
            .O(N__38892),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ));
    InMux I__8367 (
            .O(N__38889),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ));
    InMux I__8366 (
            .O(N__38886),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    InMux I__8365 (
            .O(N__38883),
            .I(N__38877));
    InMux I__8364 (
            .O(N__38882),
            .I(N__38877));
    LocalMux I__8363 (
            .O(N__38877),
            .I(N__38874));
    Span4Mux_v I__8362 (
            .O(N__38874),
            .I(N__38871));
    Odrv4 I__8361 (
            .O(N__38871),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__8360 (
            .O(N__38868),
            .I(N__38865));
    LocalMux I__8359 (
            .O(N__38865),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    CascadeMux I__8358 (
            .O(N__38862),
            .I(N__38859));
    InMux I__8357 (
            .O(N__38859),
            .I(N__38856));
    LocalMux I__8356 (
            .O(N__38856),
            .I(N__38851));
    InMux I__8355 (
            .O(N__38855),
            .I(N__38848));
    CascadeMux I__8354 (
            .O(N__38854),
            .I(N__38845));
    Span4Mux_v I__8353 (
            .O(N__38851),
            .I(N__38842));
    LocalMux I__8352 (
            .O(N__38848),
            .I(N__38839));
    InMux I__8351 (
            .O(N__38845),
            .I(N__38836));
    Span4Mux_h I__8350 (
            .O(N__38842),
            .I(N__38833));
    Span4Mux_v I__8349 (
            .O(N__38839),
            .I(N__38830));
    LocalMux I__8348 (
            .O(N__38836),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__8347 (
            .O(N__38833),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__8346 (
            .O(N__38830),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__8345 (
            .O(N__38823),
            .I(N__38819));
    InMux I__8344 (
            .O(N__38822),
            .I(N__38816));
    LocalMux I__8343 (
            .O(N__38819),
            .I(N__38813));
    LocalMux I__8342 (
            .O(N__38816),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__8341 (
            .O(N__38813),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__8340 (
            .O(N__38808),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__8339 (
            .O(N__38805),
            .I(N__38802));
    InMux I__8338 (
            .O(N__38802),
            .I(N__38799));
    LocalMux I__8337 (
            .O(N__38799),
            .I(N__38796));
    Odrv4 I__8336 (
            .O(N__38796),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ));
    InMux I__8335 (
            .O(N__38793),
            .I(N__38790));
    LocalMux I__8334 (
            .O(N__38790),
            .I(N__38786));
    InMux I__8333 (
            .O(N__38789),
            .I(N__38783));
    Span4Mux_h I__8332 (
            .O(N__38786),
            .I(N__38780));
    LocalMux I__8331 (
            .O(N__38783),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__8330 (
            .O(N__38780),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__8329 (
            .O(N__38775),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__8328 (
            .O(N__38772),
            .I(N__38768));
    InMux I__8327 (
            .O(N__38771),
            .I(N__38765));
    LocalMux I__8326 (
            .O(N__38768),
            .I(N__38762));
    LocalMux I__8325 (
            .O(N__38765),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv12 I__8324 (
            .O(N__38762),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__8323 (
            .O(N__38757),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__8322 (
            .O(N__38754),
            .I(N__38750));
    InMux I__8321 (
            .O(N__38753),
            .I(N__38747));
    LocalMux I__8320 (
            .O(N__38750),
            .I(N__38744));
    LocalMux I__8319 (
            .O(N__38747),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__8318 (
            .O(N__38744),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__8317 (
            .O(N__38739),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__8316 (
            .O(N__38736),
            .I(N__38733));
    LocalMux I__8315 (
            .O(N__38733),
            .I(N__38729));
    InMux I__8314 (
            .O(N__38732),
            .I(N__38726));
    Span4Mux_h I__8313 (
            .O(N__38729),
            .I(N__38723));
    LocalMux I__8312 (
            .O(N__38726),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__8311 (
            .O(N__38723),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__8310 (
            .O(N__38718),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    CascadeMux I__8309 (
            .O(N__38715),
            .I(N__38712));
    InMux I__8308 (
            .O(N__38712),
            .I(N__38709));
    LocalMux I__8307 (
            .O(N__38709),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__8306 (
            .O(N__38706),
            .I(N__38703));
    InMux I__8305 (
            .O(N__38703),
            .I(N__38700));
    LocalMux I__8304 (
            .O(N__38700),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    InMux I__8303 (
            .O(N__38697),
            .I(N__38694));
    LocalMux I__8302 (
            .O(N__38694),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__8301 (
            .O(N__38691),
            .I(N__38688));
    LocalMux I__8300 (
            .O(N__38688),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    CascadeMux I__8299 (
            .O(N__38685),
            .I(N__38682));
    InMux I__8298 (
            .O(N__38682),
            .I(N__38679));
    LocalMux I__8297 (
            .O(N__38679),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    InMux I__8296 (
            .O(N__38676),
            .I(N__38673));
    LocalMux I__8295 (
            .O(N__38673),
            .I(N__38670));
    Odrv12 I__8294 (
            .O(N__38670),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    CascadeMux I__8293 (
            .O(N__38667),
            .I(N__38664));
    InMux I__8292 (
            .O(N__38664),
            .I(N__38661));
    LocalMux I__8291 (
            .O(N__38661),
            .I(N__38658));
    Span4Mux_v I__8290 (
            .O(N__38658),
            .I(N__38655));
    Odrv4 I__8289 (
            .O(N__38655),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    InMux I__8288 (
            .O(N__38652),
            .I(N__38649));
    LocalMux I__8287 (
            .O(N__38649),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ));
    CascadeMux I__8286 (
            .O(N__38646),
            .I(N__38643));
    InMux I__8285 (
            .O(N__38643),
            .I(N__38640));
    LocalMux I__8284 (
            .O(N__38640),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt22 ));
    InMux I__8283 (
            .O(N__38637),
            .I(N__38634));
    LocalMux I__8282 (
            .O(N__38634),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__8281 (
            .O(N__38631),
            .I(N__38628));
    InMux I__8280 (
            .O(N__38628),
            .I(N__38625));
    LocalMux I__8279 (
            .O(N__38625),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__8278 (
            .O(N__38622),
            .I(N__38619));
    LocalMux I__8277 (
            .O(N__38619),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__8276 (
            .O(N__38616),
            .I(N__38613));
    InMux I__8275 (
            .O(N__38613),
            .I(N__38610));
    LocalMux I__8274 (
            .O(N__38610),
            .I(N__38607));
    Odrv4 I__8273 (
            .O(N__38607),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__8272 (
            .O(N__38604),
            .I(N__38601));
    InMux I__8271 (
            .O(N__38601),
            .I(N__38598));
    LocalMux I__8270 (
            .O(N__38598),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__8269 (
            .O(N__38595),
            .I(N__38592));
    LocalMux I__8268 (
            .O(N__38592),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__8267 (
            .O(N__38589),
            .I(N__38586));
    InMux I__8266 (
            .O(N__38586),
            .I(N__38583));
    LocalMux I__8265 (
            .O(N__38583),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__8264 (
            .O(N__38580),
            .I(N__38577));
    LocalMux I__8263 (
            .O(N__38577),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__8262 (
            .O(N__38574),
            .I(N__38571));
    InMux I__8261 (
            .O(N__38571),
            .I(N__38568));
    LocalMux I__8260 (
            .O(N__38568),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__8259 (
            .O(N__38565),
            .I(N__38562));
    LocalMux I__8258 (
            .O(N__38562),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__8257 (
            .O(N__38559),
            .I(N__38556));
    InMux I__8256 (
            .O(N__38556),
            .I(N__38553));
    LocalMux I__8255 (
            .O(N__38553),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__8254 (
            .O(N__38550),
            .I(N__38547));
    InMux I__8253 (
            .O(N__38547),
            .I(N__38544));
    LocalMux I__8252 (
            .O(N__38544),
            .I(N__38541));
    Odrv4 I__8251 (
            .O(N__38541),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__8250 (
            .O(N__38538),
            .I(N__38535));
    LocalMux I__8249 (
            .O(N__38535),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__8248 (
            .O(N__38532),
            .I(N__38529));
    InMux I__8247 (
            .O(N__38529),
            .I(N__38526));
    LocalMux I__8246 (
            .O(N__38526),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__8245 (
            .O(N__38523),
            .I(N__38520));
    LocalMux I__8244 (
            .O(N__38520),
            .I(N__38517));
    Odrv4 I__8243 (
            .O(N__38517),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__8242 (
            .O(N__38514),
            .I(N__38511));
    InMux I__8241 (
            .O(N__38511),
            .I(N__38508));
    LocalMux I__8240 (
            .O(N__38508),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__8239 (
            .O(N__38505),
            .I(N__38502));
    LocalMux I__8238 (
            .O(N__38502),
            .I(N__38499));
    Odrv12 I__8237 (
            .O(N__38499),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__8236 (
            .O(N__38496),
            .I(N__38493));
    InMux I__8235 (
            .O(N__38493),
            .I(N__38490));
    LocalMux I__8234 (
            .O(N__38490),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__8233 (
            .O(N__38487),
            .I(N__38484));
    LocalMux I__8232 (
            .O(N__38484),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__8231 (
            .O(N__38481),
            .I(N__38478));
    InMux I__8230 (
            .O(N__38478),
            .I(N__38475));
    LocalMux I__8229 (
            .O(N__38475),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__8228 (
            .O(N__38472),
            .I(N__38469));
    InMux I__8227 (
            .O(N__38469),
            .I(N__38466));
    LocalMux I__8226 (
            .O(N__38466),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    InMux I__8225 (
            .O(N__38463),
            .I(N__38460));
    LocalMux I__8224 (
            .O(N__38460),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__8223 (
            .O(N__38457),
            .I(N__38452));
    CascadeMux I__8222 (
            .O(N__38456),
            .I(N__38449));
    InMux I__8221 (
            .O(N__38455),
            .I(N__38443));
    InMux I__8220 (
            .O(N__38452),
            .I(N__38443));
    InMux I__8219 (
            .O(N__38449),
            .I(N__38438));
    InMux I__8218 (
            .O(N__38448),
            .I(N__38438));
    LocalMux I__8217 (
            .O(N__38443),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__8216 (
            .O(N__38438),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    IoInMux I__8215 (
            .O(N__38433),
            .I(N__38430));
    LocalMux I__8214 (
            .O(N__38430),
            .I(N__38427));
    IoSpan4Mux I__8213 (
            .O(N__38427),
            .I(N__38424));
    Sp12to4 I__8212 (
            .O(N__38424),
            .I(N__38421));
    Span12Mux_s6_v I__8211 (
            .O(N__38421),
            .I(N__38418));
    Span12Mux_v I__8210 (
            .O(N__38418),
            .I(N__38414));
    InMux I__8209 (
            .O(N__38417),
            .I(N__38411));
    Odrv12 I__8208 (
            .O(N__38414),
            .I(T12_c));
    LocalMux I__8207 (
            .O(N__38411),
            .I(T12_c));
    CascadeMux I__8206 (
            .O(N__38406),
            .I(N__38403));
    InMux I__8205 (
            .O(N__38403),
            .I(N__38399));
    InMux I__8204 (
            .O(N__38402),
            .I(N__38396));
    LocalMux I__8203 (
            .O(N__38399),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    LocalMux I__8202 (
            .O(N__38396),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    CascadeMux I__8201 (
            .O(N__38391),
            .I(N__38387));
    InMux I__8200 (
            .O(N__38390),
            .I(N__38380));
    InMux I__8199 (
            .O(N__38387),
            .I(N__38380));
    InMux I__8198 (
            .O(N__38386),
            .I(N__38377));
    InMux I__8197 (
            .O(N__38385),
            .I(N__38374));
    LocalMux I__8196 (
            .O(N__38380),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__8195 (
            .O(N__38377),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__8194 (
            .O(N__38374),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    CascadeMux I__8193 (
            .O(N__38367),
            .I(N__38363));
    InMux I__8192 (
            .O(N__38366),
            .I(N__38355));
    InMux I__8191 (
            .O(N__38363),
            .I(N__38355));
    InMux I__8190 (
            .O(N__38362),
            .I(N__38352));
    InMux I__8189 (
            .O(N__38361),
            .I(N__38347));
    InMux I__8188 (
            .O(N__38360),
            .I(N__38347));
    LocalMux I__8187 (
            .O(N__38355),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__8186 (
            .O(N__38352),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__8185 (
            .O(N__38347),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    CascadeMux I__8184 (
            .O(N__38340),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__8183 (
            .O(N__38337),
            .I(N__38331));
    InMux I__8182 (
            .O(N__38336),
            .I(N__38331));
    LocalMux I__8181 (
            .O(N__38331),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__8180 (
            .O(N__38328),
            .I(N__38325));
    InMux I__8179 (
            .O(N__38325),
            .I(N__38319));
    InMux I__8178 (
            .O(N__38324),
            .I(N__38319));
    LocalMux I__8177 (
            .O(N__38319),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__8176 (
            .O(N__38316),
            .I(N__38311));
    InMux I__8175 (
            .O(N__38315),
            .I(N__38308));
    InMux I__8174 (
            .O(N__38314),
            .I(N__38305));
    LocalMux I__8173 (
            .O(N__38311),
            .I(N__38302));
    LocalMux I__8172 (
            .O(N__38308),
            .I(N__38299));
    LocalMux I__8171 (
            .O(N__38305),
            .I(N__38296));
    Odrv12 I__8170 (
            .O(N__38302),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv12 I__8169 (
            .O(N__38299),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__8168 (
            .O(N__38296),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__8167 (
            .O(N__38289),
            .I(N__38286));
    LocalMux I__8166 (
            .O(N__38286),
            .I(N__38283));
    Odrv12 I__8165 (
            .O(N__38283),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    CascadeMux I__8164 (
            .O(N__38280),
            .I(N__38277));
    InMux I__8163 (
            .O(N__38277),
            .I(N__38271));
    InMux I__8162 (
            .O(N__38276),
            .I(N__38271));
    LocalMux I__8161 (
            .O(N__38271),
            .I(N__38267));
    InMux I__8160 (
            .O(N__38270),
            .I(N__38264));
    Span4Mux_h I__8159 (
            .O(N__38267),
            .I(N__38261));
    LocalMux I__8158 (
            .O(N__38264),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__8157 (
            .O(N__38261),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__8156 (
            .O(N__38256),
            .I(N__38252));
    InMux I__8155 (
            .O(N__38255),
            .I(N__38249));
    LocalMux I__8154 (
            .O(N__38252),
            .I(N__38242));
    LocalMux I__8153 (
            .O(N__38249),
            .I(N__38242));
    InMux I__8152 (
            .O(N__38248),
            .I(N__38239));
    InMux I__8151 (
            .O(N__38247),
            .I(N__38236));
    Span4Mux_h I__8150 (
            .O(N__38242),
            .I(N__38233));
    LocalMux I__8149 (
            .O(N__38239),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__8148 (
            .O(N__38236),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__8147 (
            .O(N__38233),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__8146 (
            .O(N__38226),
            .I(N__38220));
    ClkMux I__8145 (
            .O(N__38225),
            .I(N__38220));
    GlobalMux I__8144 (
            .O(N__38220),
            .I(N__38217));
    gio2CtrlBuf I__8143 (
            .O(N__38217),
            .I(delay_tr_input_c_g));
    InMux I__8142 (
            .O(N__38214),
            .I(N__38207));
    InMux I__8141 (
            .O(N__38213),
            .I(N__38207));
    InMux I__8140 (
            .O(N__38212),
            .I(N__38204));
    LocalMux I__8139 (
            .O(N__38207),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__8138 (
            .O(N__38204),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__8137 (
            .O(N__38199),
            .I(N__38195));
    InMux I__8136 (
            .O(N__38198),
            .I(N__38192));
    LocalMux I__8135 (
            .O(N__38195),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    LocalMux I__8134 (
            .O(N__38192),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    InMux I__8133 (
            .O(N__38187),
            .I(N__38184));
    LocalMux I__8132 (
            .O(N__38184),
            .I(\phase_controller_inst2.start_timer_tr_RNO_0_0 ));
    InMux I__8131 (
            .O(N__38181),
            .I(N__38177));
    InMux I__8130 (
            .O(N__38180),
            .I(N__38174));
    LocalMux I__8129 (
            .O(N__38177),
            .I(N__38170));
    LocalMux I__8128 (
            .O(N__38174),
            .I(N__38167));
    InMux I__8127 (
            .O(N__38173),
            .I(N__38164));
    Span4Mux_h I__8126 (
            .O(N__38170),
            .I(N__38161));
    Span4Mux_v I__8125 (
            .O(N__38167),
            .I(N__38158));
    LocalMux I__8124 (
            .O(N__38164),
            .I(N__38155));
    Span4Mux_h I__8123 (
            .O(N__38161),
            .I(N__38152));
    Span4Mux_h I__8122 (
            .O(N__38158),
            .I(N__38149));
    Span12Mux_h I__8121 (
            .O(N__38155),
            .I(N__38146));
    Span4Mux_h I__8120 (
            .O(N__38152),
            .I(N__38143));
    Span4Mux_h I__8119 (
            .O(N__38149),
            .I(N__38140));
    Odrv12 I__8118 (
            .O(N__38146),
            .I(il_max_comp2_c));
    Odrv4 I__8117 (
            .O(N__38143),
            .I(il_max_comp2_c));
    Odrv4 I__8116 (
            .O(N__38140),
            .I(il_max_comp2_c));
    InMux I__8115 (
            .O(N__38133),
            .I(N__38128));
    InMux I__8114 (
            .O(N__38132),
            .I(N__38123));
    InMux I__8113 (
            .O(N__38131),
            .I(N__38123));
    LocalMux I__8112 (
            .O(N__38128),
            .I(N__38117));
    LocalMux I__8111 (
            .O(N__38123),
            .I(N__38117));
    InMux I__8110 (
            .O(N__38122),
            .I(N__38114));
    Span4Mux_h I__8109 (
            .O(N__38117),
            .I(N__38111));
    LocalMux I__8108 (
            .O(N__38114),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__8107 (
            .O(N__38111),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__8106 (
            .O(N__38106),
            .I(N__38101));
    InMux I__8105 (
            .O(N__38105),
            .I(N__38098));
    InMux I__8104 (
            .O(N__38104),
            .I(N__38095));
    LocalMux I__8103 (
            .O(N__38101),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__8102 (
            .O(N__38098),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__8101 (
            .O(N__38095),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__8100 (
            .O(N__38088),
            .I(N__38085));
    LocalMux I__8099 (
            .O(N__38085),
            .I(N__38082));
    Odrv12 I__8098 (
            .O(N__38082),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__8097 (
            .O(N__38079),
            .I(N__38076));
    LocalMux I__8096 (
            .O(N__38076),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__8095 (
            .O(N__38073),
            .I(N__38069));
    InMux I__8094 (
            .O(N__38072),
            .I(N__38064));
    InMux I__8093 (
            .O(N__38069),
            .I(N__38064));
    LocalMux I__8092 (
            .O(N__38064),
            .I(N__38060));
    InMux I__8091 (
            .O(N__38063),
            .I(N__38057));
    Span4Mux_v I__8090 (
            .O(N__38060),
            .I(N__38054));
    LocalMux I__8089 (
            .O(N__38057),
            .I(N__38051));
    Odrv4 I__8088 (
            .O(N__38054),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__8087 (
            .O(N__38051),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__8086 (
            .O(N__38046),
            .I(N__38043));
    LocalMux I__8085 (
            .O(N__38043),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__8084 (
            .O(N__38040),
            .I(N__38019));
    InMux I__8083 (
            .O(N__38039),
            .I(N__38019));
    InMux I__8082 (
            .O(N__38038),
            .I(N__38019));
    InMux I__8081 (
            .O(N__38037),
            .I(N__38019));
    InMux I__8080 (
            .O(N__38036),
            .I(N__38019));
    InMux I__8079 (
            .O(N__38035),
            .I(N__38019));
    InMux I__8078 (
            .O(N__38034),
            .I(N__38019));
    LocalMux I__8077 (
            .O(N__38019),
            .I(N__37999));
    InMux I__8076 (
            .O(N__38018),
            .I(N__37994));
    InMux I__8075 (
            .O(N__38017),
            .I(N__37994));
    InMux I__8074 (
            .O(N__38016),
            .I(N__37991));
    InMux I__8073 (
            .O(N__38015),
            .I(N__37980));
    InMux I__8072 (
            .O(N__38014),
            .I(N__37980));
    InMux I__8071 (
            .O(N__38013),
            .I(N__37980));
    InMux I__8070 (
            .O(N__38012),
            .I(N__37980));
    InMux I__8069 (
            .O(N__38011),
            .I(N__37980));
    InMux I__8068 (
            .O(N__38010),
            .I(N__37971));
    InMux I__8067 (
            .O(N__38009),
            .I(N__37971));
    InMux I__8066 (
            .O(N__38008),
            .I(N__37971));
    InMux I__8065 (
            .O(N__38007),
            .I(N__37971));
    InMux I__8064 (
            .O(N__38006),
            .I(N__37968));
    InMux I__8063 (
            .O(N__38005),
            .I(N__37965));
    InMux I__8062 (
            .O(N__38004),
            .I(N__37958));
    InMux I__8061 (
            .O(N__38003),
            .I(N__37958));
    InMux I__8060 (
            .O(N__38002),
            .I(N__37958));
    Span4Mux_v I__8059 (
            .O(N__37999),
            .I(N__37952));
    LocalMux I__8058 (
            .O(N__37994),
            .I(N__37952));
    LocalMux I__8057 (
            .O(N__37991),
            .I(N__37947));
    LocalMux I__8056 (
            .O(N__37980),
            .I(N__37947));
    LocalMux I__8055 (
            .O(N__37971),
            .I(N__37938));
    LocalMux I__8054 (
            .O(N__37968),
            .I(N__37938));
    LocalMux I__8053 (
            .O(N__37965),
            .I(N__37938));
    LocalMux I__8052 (
            .O(N__37958),
            .I(N__37938));
    InMux I__8051 (
            .O(N__37957),
            .I(N__37935));
    Span4Mux_h I__8050 (
            .O(N__37952),
            .I(N__37932));
    Span4Mux_h I__8049 (
            .O(N__37947),
            .I(N__37929));
    Span4Mux_v I__8048 (
            .O(N__37938),
            .I(N__37926));
    LocalMux I__8047 (
            .O(N__37935),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__8046 (
            .O(N__37932),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__8045 (
            .O(N__37929),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__8044 (
            .O(N__37926),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__8043 (
            .O(N__37917),
            .I(N__37912));
    InMux I__8042 (
            .O(N__37916),
            .I(N__37909));
    InMux I__8041 (
            .O(N__37915),
            .I(N__37906));
    LocalMux I__8040 (
            .O(N__37912),
            .I(N__37901));
    LocalMux I__8039 (
            .O(N__37909),
            .I(N__37901));
    LocalMux I__8038 (
            .O(N__37906),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv12 I__8037 (
            .O(N__37901),
            .I(\current_shift_inst.un4_control_input1_25 ));
    CascadeMux I__8036 (
            .O(N__37896),
            .I(N__37893));
    InMux I__8035 (
            .O(N__37893),
            .I(N__37890));
    LocalMux I__8034 (
            .O(N__37890),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__8033 (
            .O(N__37887),
            .I(N__37884));
    LocalMux I__8032 (
            .O(N__37884),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__8031 (
            .O(N__37881),
            .I(N__37878));
    InMux I__8030 (
            .O(N__37878),
            .I(N__37875));
    LocalMux I__8029 (
            .O(N__37875),
            .I(N__37870));
    InMux I__8028 (
            .O(N__37874),
            .I(N__37867));
    InMux I__8027 (
            .O(N__37873),
            .I(N__37864));
    Span4Mux_h I__8026 (
            .O(N__37870),
            .I(N__37859));
    LocalMux I__8025 (
            .O(N__37867),
            .I(N__37859));
    LocalMux I__8024 (
            .O(N__37864),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv4 I__8023 (
            .O(N__37859),
            .I(\current_shift_inst.un4_control_input1_29 ));
    CascadeMux I__8022 (
            .O(N__37854),
            .I(N__37851));
    InMux I__8021 (
            .O(N__37851),
            .I(N__37848));
    LocalMux I__8020 (
            .O(N__37848),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    CascadeMux I__8019 (
            .O(N__37845),
            .I(N__37842));
    InMux I__8018 (
            .O(N__37842),
            .I(N__37839));
    LocalMux I__8017 (
            .O(N__37839),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    CascadeMux I__8016 (
            .O(N__37836),
            .I(N__37833));
    InMux I__8015 (
            .O(N__37833),
            .I(N__37830));
    LocalMux I__8014 (
            .O(N__37830),
            .I(N__37825));
    InMux I__8013 (
            .O(N__37829),
            .I(N__37822));
    InMux I__8012 (
            .O(N__37828),
            .I(N__37819));
    Sp12to4 I__8011 (
            .O(N__37825),
            .I(N__37814));
    LocalMux I__8010 (
            .O(N__37822),
            .I(N__37814));
    LocalMux I__8009 (
            .O(N__37819),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv12 I__8008 (
            .O(N__37814),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__8007 (
            .O(N__37809),
            .I(N__37806));
    LocalMux I__8006 (
            .O(N__37806),
            .I(N__37803));
    Odrv12 I__8005 (
            .O(N__37803),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    CascadeMux I__8004 (
            .O(N__37800),
            .I(N__37797));
    InMux I__8003 (
            .O(N__37797),
            .I(N__37794));
    LocalMux I__8002 (
            .O(N__37794),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    CascadeMux I__8001 (
            .O(N__37791),
            .I(N__37788));
    InMux I__8000 (
            .O(N__37788),
            .I(N__37785));
    LocalMux I__7999 (
            .O(N__37785),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    CascadeMux I__7998 (
            .O(N__37782),
            .I(N__37779));
    InMux I__7997 (
            .O(N__37779),
            .I(N__37776));
    LocalMux I__7996 (
            .O(N__37776),
            .I(N__37771));
    InMux I__7995 (
            .O(N__37775),
            .I(N__37768));
    InMux I__7994 (
            .O(N__37774),
            .I(N__37765));
    Span4Mux_v I__7993 (
            .O(N__37771),
            .I(N__37762));
    LocalMux I__7992 (
            .O(N__37768),
            .I(N__37759));
    LocalMux I__7991 (
            .O(N__37765),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__7990 (
            .O(N__37762),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv12 I__7989 (
            .O(N__37759),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__7988 (
            .O(N__37752),
            .I(N__37749));
    InMux I__7987 (
            .O(N__37749),
            .I(N__37746));
    LocalMux I__7986 (
            .O(N__37746),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__7985 (
            .O(N__37743),
            .I(N__37738));
    InMux I__7984 (
            .O(N__37742),
            .I(N__37735));
    InMux I__7983 (
            .O(N__37741),
            .I(N__37730));
    InMux I__7982 (
            .O(N__37738),
            .I(N__37730));
    LocalMux I__7981 (
            .O(N__37735),
            .I(N__37727));
    LocalMux I__7980 (
            .O(N__37730),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__7979 (
            .O(N__37727),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__7978 (
            .O(N__37722),
            .I(N__37719));
    LocalMux I__7977 (
            .O(N__37719),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__7976 (
            .O(N__37716),
            .I(N__37713));
    LocalMux I__7975 (
            .O(N__37713),
            .I(N__37709));
    InMux I__7974 (
            .O(N__37712),
            .I(N__37705));
    Span4Mux_v I__7973 (
            .O(N__37709),
            .I(N__37702));
    InMux I__7972 (
            .O(N__37708),
            .I(N__37699));
    LocalMux I__7971 (
            .O(N__37705),
            .I(N__37696));
    Odrv4 I__7970 (
            .O(N__37702),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__7969 (
            .O(N__37699),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv12 I__7968 (
            .O(N__37696),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__7967 (
            .O(N__37689),
            .I(N__37686));
    LocalMux I__7966 (
            .O(N__37686),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    InMux I__7965 (
            .O(N__37683),
            .I(N__37678));
    InMux I__7964 (
            .O(N__37682),
            .I(N__37675));
    InMux I__7963 (
            .O(N__37681),
            .I(N__37672));
    LocalMux I__7962 (
            .O(N__37678),
            .I(N__37669));
    LocalMux I__7961 (
            .O(N__37675),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__7960 (
            .O(N__37672),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__7959 (
            .O(N__37669),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__7958 (
            .O(N__37662),
            .I(N__37659));
    LocalMux I__7957 (
            .O(N__37659),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    CascadeMux I__7956 (
            .O(N__37656),
            .I(N__37651));
    InMux I__7955 (
            .O(N__37655),
            .I(N__37648));
    InMux I__7954 (
            .O(N__37654),
            .I(N__37645));
    InMux I__7953 (
            .O(N__37651),
            .I(N__37642));
    LocalMux I__7952 (
            .O(N__37648),
            .I(N__37639));
    LocalMux I__7951 (
            .O(N__37645),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__7950 (
            .O(N__37642),
            .I(\current_shift_inst.un4_control_input1_21 ));
    Odrv4 I__7949 (
            .O(N__37639),
            .I(\current_shift_inst.un4_control_input1_21 ));
    CascadeMux I__7948 (
            .O(N__37632),
            .I(N__37629));
    InMux I__7947 (
            .O(N__37629),
            .I(N__37626));
    LocalMux I__7946 (
            .O(N__37626),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    CascadeMux I__7945 (
            .O(N__37623),
            .I(N__37620));
    InMux I__7944 (
            .O(N__37620),
            .I(N__37617));
    LocalMux I__7943 (
            .O(N__37617),
            .I(N__37612));
    InMux I__7942 (
            .O(N__37616),
            .I(N__37609));
    InMux I__7941 (
            .O(N__37615),
            .I(N__37606));
    Span4Mux_v I__7940 (
            .O(N__37612),
            .I(N__37603));
    LocalMux I__7939 (
            .O(N__37609),
            .I(N__37600));
    LocalMux I__7938 (
            .O(N__37606),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__7937 (
            .O(N__37603),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv12 I__7936 (
            .O(N__37600),
            .I(\current_shift_inst.un4_control_input1_19 ));
    CascadeMux I__7935 (
            .O(N__37593),
            .I(N__37590));
    InMux I__7934 (
            .O(N__37590),
            .I(N__37587));
    LocalMux I__7933 (
            .O(N__37587),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    CascadeMux I__7932 (
            .O(N__37584),
            .I(N__37581));
    InMux I__7931 (
            .O(N__37581),
            .I(N__37578));
    LocalMux I__7930 (
            .O(N__37578),
            .I(N__37575));
    Span4Mux_h I__7929 (
            .O(N__37575),
            .I(N__37570));
    InMux I__7928 (
            .O(N__37574),
            .I(N__37567));
    InMux I__7927 (
            .O(N__37573),
            .I(N__37564));
    Sp12to4 I__7926 (
            .O(N__37570),
            .I(N__37559));
    LocalMux I__7925 (
            .O(N__37567),
            .I(N__37559));
    LocalMux I__7924 (
            .O(N__37564),
            .I(\current_shift_inst.un4_control_input1_9 ));
    Odrv12 I__7923 (
            .O(N__37559),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__7922 (
            .O(N__37554),
            .I(N__37551));
    LocalMux I__7921 (
            .O(N__37551),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    CascadeMux I__7920 (
            .O(N__37548),
            .I(N__37544));
    InMux I__7919 (
            .O(N__37547),
            .I(N__37541));
    InMux I__7918 (
            .O(N__37544),
            .I(N__37538));
    LocalMux I__7917 (
            .O(N__37541),
            .I(N__37532));
    LocalMux I__7916 (
            .O(N__37538),
            .I(N__37532));
    InMux I__7915 (
            .O(N__37537),
            .I(N__37529));
    Span4Mux_h I__7914 (
            .O(N__37532),
            .I(N__37526));
    LocalMux I__7913 (
            .O(N__37529),
            .I(N__37523));
    Span4Mux_h I__7912 (
            .O(N__37526),
            .I(N__37518));
    Span4Mux_v I__7911 (
            .O(N__37523),
            .I(N__37518));
    Odrv4 I__7910 (
            .O(N__37518),
            .I(\current_shift_inst.un4_control_input1_6 ));
    CascadeMux I__7909 (
            .O(N__37515),
            .I(N__37512));
    InMux I__7908 (
            .O(N__37512),
            .I(N__37509));
    LocalMux I__7907 (
            .O(N__37509),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__7906 (
            .O(N__37506),
            .I(N__37503));
    LocalMux I__7905 (
            .O(N__37503),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    CascadeMux I__7904 (
            .O(N__37500),
            .I(N__37495));
    InMux I__7903 (
            .O(N__37499),
            .I(N__37492));
    InMux I__7902 (
            .O(N__37498),
            .I(N__37487));
    InMux I__7901 (
            .O(N__37495),
            .I(N__37487));
    LocalMux I__7900 (
            .O(N__37492),
            .I(N__37484));
    LocalMux I__7899 (
            .O(N__37487),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__7898 (
            .O(N__37484),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__7897 (
            .O(N__37479),
            .I(N__37476));
    LocalMux I__7896 (
            .O(N__37476),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__7895 (
            .O(N__37473),
            .I(N__37468));
    InMux I__7894 (
            .O(N__37472),
            .I(N__37465));
    InMux I__7893 (
            .O(N__37471),
            .I(N__37462));
    LocalMux I__7892 (
            .O(N__37468),
            .I(N__37457));
    LocalMux I__7891 (
            .O(N__37465),
            .I(N__37457));
    LocalMux I__7890 (
            .O(N__37462),
            .I(N__37454));
    Span4Mux_v I__7889 (
            .O(N__37457),
            .I(N__37451));
    Span4Mux_v I__7888 (
            .O(N__37454),
            .I(N__37448));
    Odrv4 I__7887 (
            .O(N__37451),
            .I(\current_shift_inst.un4_control_input1_2 ));
    Odrv4 I__7886 (
            .O(N__37448),
            .I(\current_shift_inst.un4_control_input1_2 ));
    CascadeMux I__7885 (
            .O(N__37443),
            .I(N__37440));
    InMux I__7884 (
            .O(N__37440),
            .I(N__37437));
    LocalMux I__7883 (
            .O(N__37437),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__7882 (
            .O(N__37434),
            .I(N__37431));
    LocalMux I__7881 (
            .O(N__37431),
            .I(N__37427));
    InMux I__7880 (
            .O(N__37430),
            .I(N__37424));
    Span4Mux_h I__7879 (
            .O(N__37427),
            .I(N__37418));
    LocalMux I__7878 (
            .O(N__37424),
            .I(N__37418));
    InMux I__7877 (
            .O(N__37423),
            .I(N__37415));
    Span4Mux_v I__7876 (
            .O(N__37418),
            .I(N__37412));
    LocalMux I__7875 (
            .O(N__37415),
            .I(N__37409));
    Odrv4 I__7874 (
            .O(N__37412),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__7873 (
            .O(N__37409),
            .I(\current_shift_inst.un4_control_input1_12 ));
    CascadeMux I__7872 (
            .O(N__37404),
            .I(N__37401));
    InMux I__7871 (
            .O(N__37401),
            .I(N__37398));
    LocalMux I__7870 (
            .O(N__37398),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    CascadeMux I__7869 (
            .O(N__37395),
            .I(N__37392));
    InMux I__7868 (
            .O(N__37392),
            .I(N__37389));
    LocalMux I__7867 (
            .O(N__37389),
            .I(N__37386));
    Span4Mux_h I__7866 (
            .O(N__37386),
            .I(N__37383));
    Odrv4 I__7865 (
            .O(N__37383),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__7864 (
            .O(N__37380),
            .I(N__37376));
    InMux I__7863 (
            .O(N__37379),
            .I(N__37373));
    LocalMux I__7862 (
            .O(N__37376),
            .I(N__37369));
    LocalMux I__7861 (
            .O(N__37373),
            .I(N__37366));
    InMux I__7860 (
            .O(N__37372),
            .I(N__37363));
    Span4Mux_v I__7859 (
            .O(N__37369),
            .I(N__37360));
    Span4Mux_h I__7858 (
            .O(N__37366),
            .I(N__37357));
    LocalMux I__7857 (
            .O(N__37363),
            .I(N__37354));
    Odrv4 I__7856 (
            .O(N__37360),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__7855 (
            .O(N__37357),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__7854 (
            .O(N__37354),
            .I(\current_shift_inst.un4_control_input1_16 ));
    CascadeMux I__7853 (
            .O(N__37347),
            .I(N__37344));
    InMux I__7852 (
            .O(N__37344),
            .I(N__37341));
    LocalMux I__7851 (
            .O(N__37341),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__7850 (
            .O(N__37338),
            .I(N__37335));
    InMux I__7849 (
            .O(N__37335),
            .I(N__37332));
    LocalMux I__7848 (
            .O(N__37332),
            .I(N__37329));
    Span4Mux_h I__7847 (
            .O(N__37329),
            .I(N__37326));
    Odrv4 I__7846 (
            .O(N__37326),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    CascadeMux I__7845 (
            .O(N__37323),
            .I(N__37320));
    InMux I__7844 (
            .O(N__37320),
            .I(N__37317));
    LocalMux I__7843 (
            .O(N__37317),
            .I(N__37314));
    Span4Mux_h I__7842 (
            .O(N__37314),
            .I(N__37311));
    Odrv4 I__7841 (
            .O(N__37311),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__7840 (
            .O(N__37308),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__7839 (
            .O(N__37305),
            .I(bfn_15_16_0_));
    InMux I__7838 (
            .O(N__37302),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__7837 (
            .O(N__37299),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__7836 (
            .O(N__37296),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__7835 (
            .O(N__37293),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__7834 (
            .O(N__37290),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__7833 (
            .O(N__37287),
            .I(N__37284));
    InMux I__7832 (
            .O(N__37284),
            .I(N__37281));
    LocalMux I__7831 (
            .O(N__37281),
            .I(N__37278));
    Span4Mux_h I__7830 (
            .O(N__37278),
            .I(N__37275));
    Odrv4 I__7829 (
            .O(N__37275),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    CascadeMux I__7828 (
            .O(N__37272),
            .I(N__37269));
    InMux I__7827 (
            .O(N__37269),
            .I(N__37266));
    LocalMux I__7826 (
            .O(N__37266),
            .I(N__37263));
    Span4Mux_h I__7825 (
            .O(N__37263),
            .I(N__37260));
    Odrv4 I__7824 (
            .O(N__37260),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__7823 (
            .O(N__37257),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__7822 (
            .O(N__37254),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__7821 (
            .O(N__37251),
            .I(bfn_15_15_0_));
    InMux I__7820 (
            .O(N__37248),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__7819 (
            .O(N__37245),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__7818 (
            .O(N__37242),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    CascadeMux I__7817 (
            .O(N__37239),
            .I(N__37236));
    InMux I__7816 (
            .O(N__37236),
            .I(N__37229));
    InMux I__7815 (
            .O(N__37235),
            .I(N__37229));
    InMux I__7814 (
            .O(N__37234),
            .I(N__37226));
    LocalMux I__7813 (
            .O(N__37229),
            .I(N__37223));
    LocalMux I__7812 (
            .O(N__37226),
            .I(N__37220));
    Span4Mux_v I__7811 (
            .O(N__37223),
            .I(N__37217));
    Odrv4 I__7810 (
            .O(N__37220),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__7809 (
            .O(N__37217),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__7808 (
            .O(N__37212),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__7807 (
            .O(N__37209),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__7806 (
            .O(N__37206),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__7805 (
            .O(N__37203),
            .I(N__37200));
    LocalMux I__7804 (
            .O(N__37200),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__7803 (
            .O(N__37197),
            .I(N__37193));
    InMux I__7802 (
            .O(N__37196),
            .I(N__37190));
    LocalMux I__7801 (
            .O(N__37193),
            .I(N__37187));
    LocalMux I__7800 (
            .O(N__37190),
            .I(N__37184));
    Span4Mux_v I__7799 (
            .O(N__37187),
            .I(N__37180));
    Span4Mux_h I__7798 (
            .O(N__37184),
            .I(N__37177));
    InMux I__7797 (
            .O(N__37183),
            .I(N__37174));
    Odrv4 I__7796 (
            .O(N__37180),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__7795 (
            .O(N__37177),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__7794 (
            .O(N__37174),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__7793 (
            .O(N__37167),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__7792 (
            .O(N__37164),
            .I(N__37160));
    InMux I__7791 (
            .O(N__37163),
            .I(N__37157));
    LocalMux I__7790 (
            .O(N__37160),
            .I(N__37152));
    LocalMux I__7789 (
            .O(N__37157),
            .I(N__37152));
    Span4Mux_h I__7788 (
            .O(N__37152),
            .I(N__37148));
    InMux I__7787 (
            .O(N__37151),
            .I(N__37145));
    Odrv4 I__7786 (
            .O(N__37148),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__7785 (
            .O(N__37145),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__7784 (
            .O(N__37140),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__7783 (
            .O(N__37137),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__7782 (
            .O(N__37134),
            .I(N__37131));
    LocalMux I__7781 (
            .O(N__37131),
            .I(N__37127));
    InMux I__7780 (
            .O(N__37130),
            .I(N__37124));
    Span4Mux_h I__7779 (
            .O(N__37127),
            .I(N__37119));
    LocalMux I__7778 (
            .O(N__37124),
            .I(N__37119));
    Span4Mux_v I__7777 (
            .O(N__37119),
            .I(N__37115));
    InMux I__7776 (
            .O(N__37118),
            .I(N__37112));
    Odrv4 I__7775 (
            .O(N__37115),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__7774 (
            .O(N__37112),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__7773 (
            .O(N__37107),
            .I(bfn_15_14_0_));
    InMux I__7772 (
            .O(N__37104),
            .I(N__37101));
    LocalMux I__7771 (
            .O(N__37101),
            .I(N__37097));
    CascadeMux I__7770 (
            .O(N__37100),
            .I(N__37094));
    Span4Mux_v I__7769 (
            .O(N__37097),
            .I(N__37090));
    InMux I__7768 (
            .O(N__37094),
            .I(N__37085));
    InMux I__7767 (
            .O(N__37093),
            .I(N__37085));
    Odrv4 I__7766 (
            .O(N__37090),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__7765 (
            .O(N__37085),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__7764 (
            .O(N__37080),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__7763 (
            .O(N__37077),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    CascadeMux I__7762 (
            .O(N__37074),
            .I(N__37071));
    InMux I__7761 (
            .O(N__37071),
            .I(N__37068));
    LocalMux I__7760 (
            .O(N__37068),
            .I(N__37064));
    InMux I__7759 (
            .O(N__37067),
            .I(N__37061));
    Span4Mux_h I__7758 (
            .O(N__37064),
            .I(N__37058));
    LocalMux I__7757 (
            .O(N__37061),
            .I(N__37055));
    Span4Mux_v I__7756 (
            .O(N__37058),
            .I(N__37049));
    Span4Mux_v I__7755 (
            .O(N__37055),
            .I(N__37049));
    InMux I__7754 (
            .O(N__37054),
            .I(N__37046));
    Odrv4 I__7753 (
            .O(N__37049),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__7752 (
            .O(N__37046),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__7751 (
            .O(N__37041),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    CascadeMux I__7750 (
            .O(N__37038),
            .I(N__37035));
    InMux I__7749 (
            .O(N__37035),
            .I(N__37031));
    CascadeMux I__7748 (
            .O(N__37034),
            .I(N__37028));
    LocalMux I__7747 (
            .O(N__37031),
            .I(N__37025));
    InMux I__7746 (
            .O(N__37028),
            .I(N__37022));
    Span4Mux_v I__7745 (
            .O(N__37025),
            .I(N__37019));
    LocalMux I__7744 (
            .O(N__37022),
            .I(N__37016));
    Span4Mux_h I__7743 (
            .O(N__37019),
            .I(N__37012));
    Span4Mux_h I__7742 (
            .O(N__37016),
            .I(N__37009));
    InMux I__7741 (
            .O(N__37015),
            .I(N__37006));
    Odrv4 I__7740 (
            .O(N__37012),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__7739 (
            .O(N__37009),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__7738 (
            .O(N__37006),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__7737 (
            .O(N__36999),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__7736 (
            .O(N__36996),
            .I(N__36993));
    LocalMux I__7735 (
            .O(N__36993),
            .I(N__36990));
    Odrv4 I__7734 (
            .O(N__36990),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__7733 (
            .O(N__36987),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    CascadeMux I__7732 (
            .O(N__36984),
            .I(N__36980));
    InMux I__7731 (
            .O(N__36983),
            .I(N__36977));
    InMux I__7730 (
            .O(N__36980),
            .I(N__36974));
    LocalMux I__7729 (
            .O(N__36977),
            .I(N__36971));
    LocalMux I__7728 (
            .O(N__36974),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    Odrv4 I__7727 (
            .O(N__36971),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    CascadeMux I__7726 (
            .O(N__36966),
            .I(N__36963));
    InMux I__7725 (
            .O(N__36963),
            .I(N__36960));
    LocalMux I__7724 (
            .O(N__36960),
            .I(N__36957));
    Odrv4 I__7723 (
            .O(N__36957),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df30 ));
    InMux I__7722 (
            .O(N__36954),
            .I(N__36951));
    LocalMux I__7721 (
            .O(N__36951),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ));
    CascadeMux I__7720 (
            .O(N__36948),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__7719 (
            .O(N__36945),
            .I(N__36942));
    LocalMux I__7718 (
            .O(N__36942),
            .I(N__36939));
    Span4Mux_h I__7717 (
            .O(N__36939),
            .I(N__36936));
    Span4Mux_v I__7716 (
            .O(N__36936),
            .I(N__36932));
    InMux I__7715 (
            .O(N__36935),
            .I(N__36929));
    Odrv4 I__7714 (
            .O(N__36932),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__7713 (
            .O(N__36929),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    InMux I__7712 (
            .O(N__36924),
            .I(N__36921));
    LocalMux I__7711 (
            .O(N__36921),
            .I(N__36917));
    CascadeMux I__7710 (
            .O(N__36920),
            .I(N__36913));
    Span4Mux_v I__7709 (
            .O(N__36917),
            .I(N__36909));
    InMux I__7708 (
            .O(N__36916),
            .I(N__36906));
    InMux I__7707 (
            .O(N__36913),
            .I(N__36903));
    InMux I__7706 (
            .O(N__36912),
            .I(N__36900));
    Span4Mux_v I__7705 (
            .O(N__36909),
            .I(N__36897));
    LocalMux I__7704 (
            .O(N__36906),
            .I(N__36892));
    LocalMux I__7703 (
            .O(N__36903),
            .I(N__36892));
    LocalMux I__7702 (
            .O(N__36900),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__7701 (
            .O(N__36897),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__7700 (
            .O(N__36892),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__7699 (
            .O(N__36885),
            .I(N__36882));
    LocalMux I__7698 (
            .O(N__36882),
            .I(N__36878));
    InMux I__7697 (
            .O(N__36881),
            .I(N__36875));
    Span4Mux_v I__7696 (
            .O(N__36878),
            .I(N__36872));
    LocalMux I__7695 (
            .O(N__36875),
            .I(N__36869));
    Span4Mux_h I__7694 (
            .O(N__36872),
            .I(N__36865));
    Span4Mux_v I__7693 (
            .O(N__36869),
            .I(N__36862));
    InMux I__7692 (
            .O(N__36868),
            .I(N__36859));
    Odrv4 I__7691 (
            .O(N__36865),
            .I(\current_shift_inst.un4_control_input1_3 ));
    Odrv4 I__7690 (
            .O(N__36862),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__7689 (
            .O(N__36859),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__7688 (
            .O(N__36852),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__7687 (
            .O(N__36849),
            .I(N__36844));
    InMux I__7686 (
            .O(N__36848),
            .I(N__36841));
    InMux I__7685 (
            .O(N__36847),
            .I(N__36838));
    LocalMux I__7684 (
            .O(N__36844),
            .I(N__36833));
    LocalMux I__7683 (
            .O(N__36841),
            .I(N__36833));
    LocalMux I__7682 (
            .O(N__36838),
            .I(N__36830));
    Span4Mux_v I__7681 (
            .O(N__36833),
            .I(N__36827));
    Span4Mux_h I__7680 (
            .O(N__36830),
            .I(N__36824));
    Odrv4 I__7679 (
            .O(N__36827),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__7678 (
            .O(N__36824),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__7677 (
            .O(N__36819),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__7676 (
            .O(N__36816),
            .I(N__36811));
    InMux I__7675 (
            .O(N__36815),
            .I(N__36808));
    InMux I__7674 (
            .O(N__36814),
            .I(N__36805));
    LocalMux I__7673 (
            .O(N__36811),
            .I(N__36802));
    LocalMux I__7672 (
            .O(N__36808),
            .I(N__36797));
    LocalMux I__7671 (
            .O(N__36805),
            .I(N__36797));
    Span4Mux_h I__7670 (
            .O(N__36802),
            .I(N__36794));
    Span4Mux_v I__7669 (
            .O(N__36797),
            .I(N__36791));
    Odrv4 I__7668 (
            .O(N__36794),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__7667 (
            .O(N__36791),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__7666 (
            .O(N__36786),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__7665 (
            .O(N__36783),
            .I(N__36780));
    LocalMux I__7664 (
            .O(N__36780),
            .I(N__36777));
    Span4Mux_h I__7663 (
            .O(N__36777),
            .I(N__36774));
    Span4Mux_h I__7662 (
            .O(N__36774),
            .I(N__36771));
    Odrv4 I__7661 (
            .O(N__36771),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__7660 (
            .O(N__36768),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    CascadeMux I__7659 (
            .O(N__36765),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_));
    InMux I__7658 (
            .O(N__36762),
            .I(N__36759));
    LocalMux I__7657 (
            .O(N__36759),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__7656 (
            .O(N__36756),
            .I(N__36753));
    LocalMux I__7655 (
            .O(N__36753),
            .I(N__36749));
    InMux I__7654 (
            .O(N__36752),
            .I(N__36746));
    Odrv4 I__7653 (
            .O(N__36749),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    LocalMux I__7652 (
            .O(N__36746),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    CascadeMux I__7651 (
            .O(N__36741),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17_cascade_));
    InMux I__7650 (
            .O(N__36738),
            .I(N__36730));
    InMux I__7649 (
            .O(N__36737),
            .I(N__36730));
    InMux I__7648 (
            .O(N__36736),
            .I(N__36727));
    InMux I__7647 (
            .O(N__36735),
            .I(N__36724));
    LocalMux I__7646 (
            .O(N__36730),
            .I(N__36719));
    LocalMux I__7645 (
            .O(N__36727),
            .I(N__36719));
    LocalMux I__7644 (
            .O(N__36724),
            .I(N__36716));
    Span4Mux_v I__7643 (
            .O(N__36719),
            .I(N__36713));
    Odrv4 I__7642 (
            .O(N__36716),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv4 I__7641 (
            .O(N__36713),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__7640 (
            .O(N__36708),
            .I(N__36705));
    LocalMux I__7639 (
            .O(N__36705),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    CascadeMux I__7638 (
            .O(N__36702),
            .I(N__36699));
    InMux I__7637 (
            .O(N__36699),
            .I(N__36693));
    InMux I__7636 (
            .O(N__36698),
            .I(N__36693));
    LocalMux I__7635 (
            .O(N__36693),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__7634 (
            .O(N__36690),
            .I(N__36687));
    InMux I__7633 (
            .O(N__36687),
            .I(N__36684));
    LocalMux I__7632 (
            .O(N__36684),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    InMux I__7631 (
            .O(N__36681),
            .I(N__36678));
    LocalMux I__7630 (
            .O(N__36678),
            .I(N__36674));
    InMux I__7629 (
            .O(N__36677),
            .I(N__36671));
    Odrv12 I__7628 (
            .O(N__36674),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    LocalMux I__7627 (
            .O(N__36671),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    CascadeMux I__7626 (
            .O(N__36666),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_));
    InMux I__7625 (
            .O(N__36663),
            .I(N__36658));
    InMux I__7624 (
            .O(N__36662),
            .I(N__36653));
    InMux I__7623 (
            .O(N__36661),
            .I(N__36653));
    LocalMux I__7622 (
            .O(N__36658),
            .I(N__36649));
    LocalMux I__7621 (
            .O(N__36653),
            .I(N__36646));
    InMux I__7620 (
            .O(N__36652),
            .I(N__36643));
    Sp12to4 I__7619 (
            .O(N__36649),
            .I(N__36640));
    Span4Mux_h I__7618 (
            .O(N__36646),
            .I(N__36637));
    LocalMux I__7617 (
            .O(N__36643),
            .I(N__36634));
    Odrv12 I__7616 (
            .O(N__36640),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv4 I__7615 (
            .O(N__36637),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv4 I__7614 (
            .O(N__36634),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__7613 (
            .O(N__36627),
            .I(N__36621));
    InMux I__7612 (
            .O(N__36626),
            .I(N__36621));
    LocalMux I__7611 (
            .O(N__36621),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__7610 (
            .O(N__36618),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12_cascade_));
    InMux I__7609 (
            .O(N__36615),
            .I(N__36612));
    LocalMux I__7608 (
            .O(N__36612),
            .I(N__36608));
    InMux I__7607 (
            .O(N__36611),
            .I(N__36605));
    Span4Mux_h I__7606 (
            .O(N__36608),
            .I(N__36599));
    LocalMux I__7605 (
            .O(N__36605),
            .I(N__36599));
    InMux I__7604 (
            .O(N__36604),
            .I(N__36596));
    Span4Mux_v I__7603 (
            .O(N__36599),
            .I(N__36593));
    LocalMux I__7602 (
            .O(N__36596),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    Odrv4 I__7601 (
            .O(N__36593),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    CascadeMux I__7600 (
            .O(N__36588),
            .I(N__36585));
    InMux I__7599 (
            .O(N__36585),
            .I(N__36582));
    LocalMux I__7598 (
            .O(N__36582),
            .I(N__36579));
    Span4Mux_v I__7597 (
            .O(N__36579),
            .I(N__36576));
    Odrv4 I__7596 (
            .O(N__36576),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt20 ));
    CascadeMux I__7595 (
            .O(N__36573),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_));
    InMux I__7594 (
            .O(N__36570),
            .I(N__36564));
    InMux I__7593 (
            .O(N__36569),
            .I(N__36564));
    LocalMux I__7592 (
            .O(N__36564),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    CascadeMux I__7591 (
            .O(N__36561),
            .I(N__36558));
    InMux I__7590 (
            .O(N__36558),
            .I(N__36552));
    InMux I__7589 (
            .O(N__36557),
            .I(N__36552));
    LocalMux I__7588 (
            .O(N__36552),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    InMux I__7587 (
            .O(N__36549),
            .I(N__36546));
    LocalMux I__7586 (
            .O(N__36546),
            .I(N__36543));
    Odrv4 I__7585 (
            .O(N__36543),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ));
    InMux I__7584 (
            .O(N__36540),
            .I(N__36536));
    InMux I__7583 (
            .O(N__36539),
            .I(N__36532));
    LocalMux I__7582 (
            .O(N__36536),
            .I(N__36529));
    InMux I__7581 (
            .O(N__36535),
            .I(N__36526));
    LocalMux I__7580 (
            .O(N__36532),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__7579 (
            .O(N__36529),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    LocalMux I__7578 (
            .O(N__36526),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__7577 (
            .O(N__36519),
            .I(N__36516));
    LocalMux I__7576 (
            .O(N__36516),
            .I(N__36510));
    InMux I__7575 (
            .O(N__36515),
            .I(N__36507));
    InMux I__7574 (
            .O(N__36514),
            .I(N__36502));
    InMux I__7573 (
            .O(N__36513),
            .I(N__36502));
    Odrv4 I__7572 (
            .O(N__36510),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__7571 (
            .O(N__36507),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__7570 (
            .O(N__36502),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__7569 (
            .O(N__36495),
            .I(N__36492));
    LocalMux I__7568 (
            .O(N__36492),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__7567 (
            .O(N__36489),
            .I(N__36485));
    InMux I__7566 (
            .O(N__36488),
            .I(N__36481));
    LocalMux I__7565 (
            .O(N__36485),
            .I(N__36478));
    InMux I__7564 (
            .O(N__36484),
            .I(N__36475));
    LocalMux I__7563 (
            .O(N__36481),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv4 I__7562 (
            .O(N__36478),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    LocalMux I__7561 (
            .O(N__36475),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__7560 (
            .O(N__36468),
            .I(N__36464));
    InMux I__7559 (
            .O(N__36467),
            .I(N__36461));
    LocalMux I__7558 (
            .O(N__36464),
            .I(N__36454));
    LocalMux I__7557 (
            .O(N__36461),
            .I(N__36454));
    InMux I__7556 (
            .O(N__36460),
            .I(N__36451));
    InMux I__7555 (
            .O(N__36459),
            .I(N__36448));
    Span4Mux_v I__7554 (
            .O(N__36454),
            .I(N__36441));
    LocalMux I__7553 (
            .O(N__36451),
            .I(N__36441));
    LocalMux I__7552 (
            .O(N__36448),
            .I(N__36441));
    Odrv4 I__7551 (
            .O(N__36441),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    CascadeMux I__7550 (
            .O(N__36438),
            .I(N__36435));
    InMux I__7549 (
            .O(N__36435),
            .I(N__36432));
    LocalMux I__7548 (
            .O(N__36432),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__7547 (
            .O(N__36429),
            .I(N__36425));
    InMux I__7546 (
            .O(N__36428),
            .I(N__36421));
    LocalMux I__7545 (
            .O(N__36425),
            .I(N__36418));
    InMux I__7544 (
            .O(N__36424),
            .I(N__36415));
    LocalMux I__7543 (
            .O(N__36421),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    Odrv4 I__7542 (
            .O(N__36418),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    LocalMux I__7541 (
            .O(N__36415),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__7540 (
            .O(N__36408),
            .I(N__36404));
    InMux I__7539 (
            .O(N__36407),
            .I(N__36401));
    LocalMux I__7538 (
            .O(N__36404),
            .I(N__36394));
    LocalMux I__7537 (
            .O(N__36401),
            .I(N__36394));
    InMux I__7536 (
            .O(N__36400),
            .I(N__36389));
    InMux I__7535 (
            .O(N__36399),
            .I(N__36389));
    Span4Mux_v I__7534 (
            .O(N__36394),
            .I(N__36384));
    LocalMux I__7533 (
            .O(N__36389),
            .I(N__36384));
    Odrv4 I__7532 (
            .O(N__36384),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__7531 (
            .O(N__36381),
            .I(N__36378));
    LocalMux I__7530 (
            .O(N__36378),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__7529 (
            .O(N__36375),
            .I(N__36372));
    InMux I__7528 (
            .O(N__36372),
            .I(N__36366));
    InMux I__7527 (
            .O(N__36371),
            .I(N__36363));
    InMux I__7526 (
            .O(N__36370),
            .I(N__36358));
    InMux I__7525 (
            .O(N__36369),
            .I(N__36358));
    LocalMux I__7524 (
            .O(N__36366),
            .I(N__36355));
    LocalMux I__7523 (
            .O(N__36363),
            .I(N__36352));
    LocalMux I__7522 (
            .O(N__36358),
            .I(N__36349));
    Span4Mux_h I__7521 (
            .O(N__36355),
            .I(N__36346));
    Odrv4 I__7520 (
            .O(N__36352),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv4 I__7519 (
            .O(N__36349),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv4 I__7518 (
            .O(N__36346),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__7517 (
            .O(N__36339),
            .I(N__36336));
    LocalMux I__7516 (
            .O(N__36336),
            .I(N__36333));
    Span4Mux_h I__7515 (
            .O(N__36333),
            .I(N__36329));
    InMux I__7514 (
            .O(N__36332),
            .I(N__36326));
    Odrv4 I__7513 (
            .O(N__36329),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__7512 (
            .O(N__36326),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    InMux I__7511 (
            .O(N__36321),
            .I(N__36315));
    InMux I__7510 (
            .O(N__36320),
            .I(N__36315));
    LocalMux I__7509 (
            .O(N__36315),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ));
    InMux I__7508 (
            .O(N__36312),
            .I(N__36309));
    LocalMux I__7507 (
            .O(N__36309),
            .I(N__36306));
    Span4Mux_v I__7506 (
            .O(N__36306),
            .I(N__36302));
    InMux I__7505 (
            .O(N__36305),
            .I(N__36299));
    Odrv4 I__7504 (
            .O(N__36302),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__7503 (
            .O(N__36299),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    InMux I__7502 (
            .O(N__36294),
            .I(N__36289));
    InMux I__7501 (
            .O(N__36293),
            .I(N__36284));
    InMux I__7500 (
            .O(N__36292),
            .I(N__36284));
    LocalMux I__7499 (
            .O(N__36289),
            .I(N__36280));
    LocalMux I__7498 (
            .O(N__36284),
            .I(N__36277));
    InMux I__7497 (
            .O(N__36283),
            .I(N__36274));
    Odrv4 I__7496 (
            .O(N__36280),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    Odrv4 I__7495 (
            .O(N__36277),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__7494 (
            .O(N__36274),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    CascadeMux I__7493 (
            .O(N__36267),
            .I(N__36264));
    InMux I__7492 (
            .O(N__36264),
            .I(N__36258));
    InMux I__7491 (
            .O(N__36263),
            .I(N__36258));
    LocalMux I__7490 (
            .O(N__36258),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ));
    InMux I__7489 (
            .O(N__36255),
            .I(N__36251));
    InMux I__7488 (
            .O(N__36254),
            .I(N__36248));
    LocalMux I__7487 (
            .O(N__36251),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__7486 (
            .O(N__36248),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    InMux I__7485 (
            .O(N__36243),
            .I(N__36240));
    LocalMux I__7484 (
            .O(N__36240),
            .I(N__36237));
    Span4Mux_v I__7483 (
            .O(N__36237),
            .I(N__36234));
    Odrv4 I__7482 (
            .O(N__36234),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__7481 (
            .O(N__36231),
            .I(N__36227));
    InMux I__7480 (
            .O(N__36230),
            .I(N__36224));
    InMux I__7479 (
            .O(N__36227),
            .I(N__36221));
    LocalMux I__7478 (
            .O(N__36224),
            .I(N__36217));
    LocalMux I__7477 (
            .O(N__36221),
            .I(N__36214));
    InMux I__7476 (
            .O(N__36220),
            .I(N__36211));
    Odrv4 I__7475 (
            .O(N__36217),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__7474 (
            .O(N__36214),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__7473 (
            .O(N__36211),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    CEMux I__7472 (
            .O(N__36204),
            .I(N__36200));
    CEMux I__7471 (
            .O(N__36203),
            .I(N__36197));
    LocalMux I__7470 (
            .O(N__36200),
            .I(N__36191));
    LocalMux I__7469 (
            .O(N__36197),
            .I(N__36188));
    CEMux I__7468 (
            .O(N__36196),
            .I(N__36185));
    CEMux I__7467 (
            .O(N__36195),
            .I(N__36182));
    CEMux I__7466 (
            .O(N__36194),
            .I(N__36179));
    Span4Mux_v I__7465 (
            .O(N__36191),
            .I(N__36175));
    Span4Mux_h I__7464 (
            .O(N__36188),
            .I(N__36172));
    LocalMux I__7463 (
            .O(N__36185),
            .I(N__36169));
    LocalMux I__7462 (
            .O(N__36182),
            .I(N__36166));
    LocalMux I__7461 (
            .O(N__36179),
            .I(N__36163));
    CEMux I__7460 (
            .O(N__36178),
            .I(N__36160));
    Span4Mux_v I__7459 (
            .O(N__36175),
            .I(N__36157));
    Span4Mux_v I__7458 (
            .O(N__36172),
            .I(N__36154));
    Span4Mux_v I__7457 (
            .O(N__36169),
            .I(N__36145));
    Span4Mux_v I__7456 (
            .O(N__36166),
            .I(N__36145));
    Span4Mux_h I__7455 (
            .O(N__36163),
            .I(N__36145));
    LocalMux I__7454 (
            .O(N__36160),
            .I(N__36145));
    Span4Mux_v I__7453 (
            .O(N__36157),
            .I(N__36142));
    Span4Mux_v I__7452 (
            .O(N__36154),
            .I(N__36139));
    Span4Mux_v I__7451 (
            .O(N__36145),
            .I(N__36136));
    Span4Mux_v I__7450 (
            .O(N__36142),
            .I(N__36133));
    Span4Mux_v I__7449 (
            .O(N__36139),
            .I(N__36130));
    Span4Mux_v I__7448 (
            .O(N__36136),
            .I(N__36127));
    Odrv4 I__7447 (
            .O(N__36133),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv4 I__7446 (
            .O(N__36130),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    Odrv4 I__7445 (
            .O(N__36127),
            .I(\delay_measurement_inst.delay_tr_timer.N_200_i ));
    InMux I__7444 (
            .O(N__36120),
            .I(N__36114));
    InMux I__7443 (
            .O(N__36119),
            .I(N__36114));
    LocalMux I__7442 (
            .O(N__36114),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__7441 (
            .O(N__36111),
            .I(N__36108));
    InMux I__7440 (
            .O(N__36108),
            .I(N__36102));
    InMux I__7439 (
            .O(N__36107),
            .I(N__36102));
    LocalMux I__7438 (
            .O(N__36102),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    InMux I__7437 (
            .O(N__36099),
            .I(N__36096));
    LocalMux I__7436 (
            .O(N__36096),
            .I(N__36093));
    Odrv4 I__7435 (
            .O(N__36093),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ));
    CascadeMux I__7434 (
            .O(N__36090),
            .I(N__36085));
    InMux I__7433 (
            .O(N__36089),
            .I(N__36082));
    InMux I__7432 (
            .O(N__36088),
            .I(N__36070));
    InMux I__7431 (
            .O(N__36085),
            .I(N__36070));
    LocalMux I__7430 (
            .O(N__36082),
            .I(N__36067));
    InMux I__7429 (
            .O(N__36081),
            .I(N__36052));
    InMux I__7428 (
            .O(N__36080),
            .I(N__36052));
    InMux I__7427 (
            .O(N__36079),
            .I(N__36052));
    InMux I__7426 (
            .O(N__36078),
            .I(N__36052));
    InMux I__7425 (
            .O(N__36077),
            .I(N__36052));
    InMux I__7424 (
            .O(N__36076),
            .I(N__36052));
    InMux I__7423 (
            .O(N__36075),
            .I(N__36052));
    LocalMux I__7422 (
            .O(N__36070),
            .I(N__36049));
    Span4Mux_h I__7421 (
            .O(N__36067),
            .I(N__36044));
    LocalMux I__7420 (
            .O(N__36052),
            .I(N__36044));
    Span4Mux_h I__7419 (
            .O(N__36049),
            .I(N__36041));
    Span4Mux_h I__7418 (
            .O(N__36044),
            .I(N__36038));
    Span4Mux_h I__7417 (
            .O(N__36041),
            .I(N__36035));
    Span4Mux_h I__7416 (
            .O(N__36038),
            .I(N__36032));
    Span4Mux_h I__7415 (
            .O(N__36035),
            .I(N__36029));
    Span4Mux_h I__7414 (
            .O(N__36032),
            .I(N__36026));
    Odrv4 I__7413 (
            .O(N__36029),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__7412 (
            .O(N__36026),
            .I(\pwm_generator_inst.N_16 ));
    InMux I__7411 (
            .O(N__36021),
            .I(N__35993));
    InMux I__7410 (
            .O(N__36020),
            .I(N__35993));
    InMux I__7409 (
            .O(N__36019),
            .I(N__35986));
    InMux I__7408 (
            .O(N__36018),
            .I(N__35986));
    InMux I__7407 (
            .O(N__36017),
            .I(N__35986));
    InMux I__7406 (
            .O(N__36016),
            .I(N__35969));
    InMux I__7405 (
            .O(N__36015),
            .I(N__35969));
    InMux I__7404 (
            .O(N__36014),
            .I(N__35969));
    InMux I__7403 (
            .O(N__36013),
            .I(N__35969));
    InMux I__7402 (
            .O(N__36012),
            .I(N__35969));
    InMux I__7401 (
            .O(N__36011),
            .I(N__35969));
    InMux I__7400 (
            .O(N__36010),
            .I(N__35969));
    InMux I__7399 (
            .O(N__36009),
            .I(N__35969));
    InMux I__7398 (
            .O(N__36008),
            .I(N__35954));
    InMux I__7397 (
            .O(N__36007),
            .I(N__35954));
    InMux I__7396 (
            .O(N__36006),
            .I(N__35954));
    InMux I__7395 (
            .O(N__36005),
            .I(N__35954));
    InMux I__7394 (
            .O(N__36004),
            .I(N__35954));
    InMux I__7393 (
            .O(N__36003),
            .I(N__35954));
    InMux I__7392 (
            .O(N__36002),
            .I(N__35954));
    CascadeMux I__7391 (
            .O(N__36001),
            .I(N__35947));
    CascadeMux I__7390 (
            .O(N__36000),
            .I(N__35944));
    CascadeMux I__7389 (
            .O(N__35999),
            .I(N__35940));
    CascadeMux I__7388 (
            .O(N__35998),
            .I(N__35936));
    LocalMux I__7387 (
            .O(N__35993),
            .I(N__35931));
    LocalMux I__7386 (
            .O(N__35986),
            .I(N__35931));
    LocalMux I__7385 (
            .O(N__35969),
            .I(N__35926));
    LocalMux I__7384 (
            .O(N__35954),
            .I(N__35926));
    InMux I__7383 (
            .O(N__35953),
            .I(N__35921));
    InMux I__7382 (
            .O(N__35952),
            .I(N__35921));
    InMux I__7381 (
            .O(N__35951),
            .I(N__35906));
    InMux I__7380 (
            .O(N__35950),
            .I(N__35906));
    InMux I__7379 (
            .O(N__35947),
            .I(N__35906));
    InMux I__7378 (
            .O(N__35944),
            .I(N__35906));
    InMux I__7377 (
            .O(N__35943),
            .I(N__35906));
    InMux I__7376 (
            .O(N__35940),
            .I(N__35906));
    InMux I__7375 (
            .O(N__35939),
            .I(N__35906));
    InMux I__7374 (
            .O(N__35936),
            .I(N__35903));
    Span4Mux_v I__7373 (
            .O(N__35931),
            .I(N__35899));
    Span4Mux_v I__7372 (
            .O(N__35926),
            .I(N__35896));
    LocalMux I__7371 (
            .O(N__35921),
            .I(N__35893));
    LocalMux I__7370 (
            .O(N__35906),
            .I(N__35888));
    LocalMux I__7369 (
            .O(N__35903),
            .I(N__35888));
    CascadeMux I__7368 (
            .O(N__35902),
            .I(N__35885));
    Span4Mux_h I__7367 (
            .O(N__35899),
            .I(N__35881));
    Sp12to4 I__7366 (
            .O(N__35896),
            .I(N__35878));
    Span4Mux_h I__7365 (
            .O(N__35893),
            .I(N__35875));
    Span4Mux_h I__7364 (
            .O(N__35888),
            .I(N__35872));
    InMux I__7363 (
            .O(N__35885),
            .I(N__35867));
    InMux I__7362 (
            .O(N__35884),
            .I(N__35867));
    Sp12to4 I__7361 (
            .O(N__35881),
            .I(N__35862));
    Span12Mux_s8_h I__7360 (
            .O(N__35878),
            .I(N__35862));
    Odrv4 I__7359 (
            .O(N__35875),
            .I(N_19_1));
    Odrv4 I__7358 (
            .O(N__35872),
            .I(N_19_1));
    LocalMux I__7357 (
            .O(N__35867),
            .I(N_19_1));
    Odrv12 I__7356 (
            .O(N__35862),
            .I(N_19_1));
    InMux I__7355 (
            .O(N__35853),
            .I(N__35847));
    InMux I__7354 (
            .O(N__35852),
            .I(N__35847));
    LocalMux I__7353 (
            .O(N__35847),
            .I(N__35843));
    InMux I__7352 (
            .O(N__35846),
            .I(N__35833));
    Span4Mux_v I__7351 (
            .O(N__35843),
            .I(N__35830));
    InMux I__7350 (
            .O(N__35842),
            .I(N__35815));
    InMux I__7349 (
            .O(N__35841),
            .I(N__35815));
    InMux I__7348 (
            .O(N__35840),
            .I(N__35815));
    InMux I__7347 (
            .O(N__35839),
            .I(N__35815));
    InMux I__7346 (
            .O(N__35838),
            .I(N__35815));
    InMux I__7345 (
            .O(N__35837),
            .I(N__35815));
    InMux I__7344 (
            .O(N__35836),
            .I(N__35815));
    LocalMux I__7343 (
            .O(N__35833),
            .I(N__35812));
    Sp12to4 I__7342 (
            .O(N__35830),
            .I(N__35805));
    LocalMux I__7341 (
            .O(N__35815),
            .I(N__35805));
    Sp12to4 I__7340 (
            .O(N__35812),
            .I(N__35805));
    Odrv12 I__7339 (
            .O(N__35805),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__7338 (
            .O(N__35802),
            .I(N__35799));
    InMux I__7337 (
            .O(N__35799),
            .I(N__35796));
    LocalMux I__7336 (
            .O(N__35796),
            .I(N__35793));
    Odrv4 I__7335 (
            .O(N__35793),
            .I(\pwm_generator_inst.threshold_0 ));
    InMux I__7334 (
            .O(N__35790),
            .I(N__35787));
    LocalMux I__7333 (
            .O(N__35787),
            .I(N__35783));
    InMux I__7332 (
            .O(N__35786),
            .I(N__35780));
    Span12Mux_h I__7331 (
            .O(N__35783),
            .I(N__35777));
    LocalMux I__7330 (
            .O(N__35780),
            .I(N__35774));
    Odrv12 I__7329 (
            .O(N__35777),
            .I(state_ns_i_a3_1));
    Odrv4 I__7328 (
            .O(N__35774),
            .I(state_ns_i_a3_1));
    IoInMux I__7327 (
            .O(N__35769),
            .I(N__35766));
    LocalMux I__7326 (
            .O(N__35766),
            .I(N__35763));
    IoSpan4Mux I__7325 (
            .O(N__35763),
            .I(N__35760));
    Span4Mux_s1_v I__7324 (
            .O(N__35760),
            .I(N__35757));
    Sp12to4 I__7323 (
            .O(N__35757),
            .I(N__35754));
    Span12Mux_v I__7322 (
            .O(N__35754),
            .I(N__35751));
    Span12Mux_v I__7321 (
            .O(N__35751),
            .I(N__35747));
    InMux I__7320 (
            .O(N__35750),
            .I(N__35744));
    Odrv12 I__7319 (
            .O(N__35747),
            .I(T45_c));
    LocalMux I__7318 (
            .O(N__35744),
            .I(T45_c));
    InMux I__7317 (
            .O(N__35739),
            .I(N__35735));
    InMux I__7316 (
            .O(N__35738),
            .I(N__35732));
    LocalMux I__7315 (
            .O(N__35735),
            .I(N__35726));
    LocalMux I__7314 (
            .O(N__35732),
            .I(N__35726));
    InMux I__7313 (
            .O(N__35731),
            .I(N__35723));
    Span4Mux_v I__7312 (
            .O(N__35726),
            .I(N__35718));
    LocalMux I__7311 (
            .O(N__35723),
            .I(N__35718));
    Span4Mux_h I__7310 (
            .O(N__35718),
            .I(N__35715));
    Span4Mux_h I__7309 (
            .O(N__35715),
            .I(N__35712));
    Odrv4 I__7308 (
            .O(N__35712),
            .I(il_min_comp2_c));
    InMux I__7307 (
            .O(N__35709),
            .I(N__35705));
    InMux I__7306 (
            .O(N__35708),
            .I(N__35702));
    LocalMux I__7305 (
            .O(N__35705),
            .I(N__35699));
    LocalMux I__7304 (
            .O(N__35702),
            .I(N__35696));
    Span4Mux_v I__7303 (
            .O(N__35699),
            .I(N__35691));
    Span4Mux_v I__7302 (
            .O(N__35696),
            .I(N__35691));
    Odrv4 I__7301 (
            .O(N__35691),
            .I(\phase_controller_inst2.time_passed_RNIG7JF ));
    InMux I__7300 (
            .O(N__35688),
            .I(N__35685));
    LocalMux I__7299 (
            .O(N__35685),
            .I(N__35682));
    Span4Mux_v I__7298 (
            .O(N__35682),
            .I(N__35679));
    Odrv4 I__7297 (
            .O(N__35679),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__7296 (
            .O(N__35676),
            .I(N__35672));
    InMux I__7295 (
            .O(N__35675),
            .I(N__35665));
    LocalMux I__7294 (
            .O(N__35672),
            .I(N__35654));
    InMux I__7293 (
            .O(N__35671),
            .I(N__35651));
    InMux I__7292 (
            .O(N__35670),
            .I(N__35646));
    InMux I__7291 (
            .O(N__35669),
            .I(N__35646));
    InMux I__7290 (
            .O(N__35668),
            .I(N__35643));
    LocalMux I__7289 (
            .O(N__35665),
            .I(N__35637));
    InMux I__7288 (
            .O(N__35664),
            .I(N__35634));
    InMux I__7287 (
            .O(N__35663),
            .I(N__35627));
    InMux I__7286 (
            .O(N__35662),
            .I(N__35627));
    InMux I__7285 (
            .O(N__35661),
            .I(N__35627));
    InMux I__7284 (
            .O(N__35660),
            .I(N__35618));
    InMux I__7283 (
            .O(N__35659),
            .I(N__35618));
    InMux I__7282 (
            .O(N__35658),
            .I(N__35618));
    InMux I__7281 (
            .O(N__35657),
            .I(N__35618));
    Span4Mux_v I__7280 (
            .O(N__35654),
            .I(N__35611));
    LocalMux I__7279 (
            .O(N__35651),
            .I(N__35611));
    LocalMux I__7278 (
            .O(N__35646),
            .I(N__35611));
    LocalMux I__7277 (
            .O(N__35643),
            .I(N__35608));
    InMux I__7276 (
            .O(N__35642),
            .I(N__35604));
    InMux I__7275 (
            .O(N__35641),
            .I(N__35601));
    InMux I__7274 (
            .O(N__35640),
            .I(N__35598));
    Span4Mux_v I__7273 (
            .O(N__35637),
            .I(N__35572));
    LocalMux I__7272 (
            .O(N__35634),
            .I(N__35572));
    LocalMux I__7271 (
            .O(N__35627),
            .I(N__35572));
    LocalMux I__7270 (
            .O(N__35618),
            .I(N__35572));
    Span4Mux_v I__7269 (
            .O(N__35611),
            .I(N__35569));
    Span4Mux_v I__7268 (
            .O(N__35608),
            .I(N__35566));
    InMux I__7267 (
            .O(N__35607),
            .I(N__35563));
    LocalMux I__7266 (
            .O(N__35604),
            .I(N__35560));
    LocalMux I__7265 (
            .O(N__35601),
            .I(N__35555));
    LocalMux I__7264 (
            .O(N__35598),
            .I(N__35555));
    InMux I__7263 (
            .O(N__35597),
            .I(N__35548));
    InMux I__7262 (
            .O(N__35596),
            .I(N__35548));
    InMux I__7261 (
            .O(N__35595),
            .I(N__35548));
    InMux I__7260 (
            .O(N__35594),
            .I(N__35539));
    InMux I__7259 (
            .O(N__35593),
            .I(N__35539));
    InMux I__7258 (
            .O(N__35592),
            .I(N__35539));
    InMux I__7257 (
            .O(N__35591),
            .I(N__35539));
    CascadeMux I__7256 (
            .O(N__35590),
            .I(N__35534));
    CascadeMux I__7255 (
            .O(N__35589),
            .I(N__35530));
    CascadeMux I__7254 (
            .O(N__35588),
            .I(N__35526));
    CascadeMux I__7253 (
            .O(N__35587),
            .I(N__35521));
    CascadeMux I__7252 (
            .O(N__35586),
            .I(N__35517));
    CascadeMux I__7251 (
            .O(N__35585),
            .I(N__35513));
    CascadeMux I__7250 (
            .O(N__35584),
            .I(N__35509));
    InMux I__7249 (
            .O(N__35583),
            .I(N__35495));
    InMux I__7248 (
            .O(N__35582),
            .I(N__35495));
    InMux I__7247 (
            .O(N__35581),
            .I(N__35492));
    Span4Mux_v I__7246 (
            .O(N__35572),
            .I(N__35489));
    Span4Mux_v I__7245 (
            .O(N__35569),
            .I(N__35484));
    Span4Mux_v I__7244 (
            .O(N__35566),
            .I(N__35484));
    LocalMux I__7243 (
            .O(N__35563),
            .I(N__35481));
    Span4Mux_v I__7242 (
            .O(N__35560),
            .I(N__35472));
    Span4Mux_v I__7241 (
            .O(N__35555),
            .I(N__35472));
    LocalMux I__7240 (
            .O(N__35548),
            .I(N__35472));
    LocalMux I__7239 (
            .O(N__35539),
            .I(N__35472));
    CascadeMux I__7238 (
            .O(N__35538),
            .I(N__35468));
    InMux I__7237 (
            .O(N__35537),
            .I(N__35452));
    InMux I__7236 (
            .O(N__35534),
            .I(N__35452));
    InMux I__7235 (
            .O(N__35533),
            .I(N__35452));
    InMux I__7234 (
            .O(N__35530),
            .I(N__35452));
    InMux I__7233 (
            .O(N__35529),
            .I(N__35452));
    InMux I__7232 (
            .O(N__35526),
            .I(N__35452));
    InMux I__7231 (
            .O(N__35525),
            .I(N__35452));
    InMux I__7230 (
            .O(N__35524),
            .I(N__35435));
    InMux I__7229 (
            .O(N__35521),
            .I(N__35435));
    InMux I__7228 (
            .O(N__35520),
            .I(N__35435));
    InMux I__7227 (
            .O(N__35517),
            .I(N__35435));
    InMux I__7226 (
            .O(N__35516),
            .I(N__35435));
    InMux I__7225 (
            .O(N__35513),
            .I(N__35435));
    InMux I__7224 (
            .O(N__35512),
            .I(N__35435));
    InMux I__7223 (
            .O(N__35509),
            .I(N__35435));
    InMux I__7222 (
            .O(N__35508),
            .I(N__35430));
    InMux I__7221 (
            .O(N__35507),
            .I(N__35430));
    CascadeMux I__7220 (
            .O(N__35506),
            .I(N__35427));
    CascadeMux I__7219 (
            .O(N__35505),
            .I(N__35423));
    CascadeMux I__7218 (
            .O(N__35504),
            .I(N__35419));
    CascadeMux I__7217 (
            .O(N__35503),
            .I(N__35415));
    CascadeMux I__7216 (
            .O(N__35502),
            .I(N__35410));
    CascadeMux I__7215 (
            .O(N__35501),
            .I(N__35406));
    CascadeMux I__7214 (
            .O(N__35500),
            .I(N__35402));
    LocalMux I__7213 (
            .O(N__35495),
            .I(N__35396));
    LocalMux I__7212 (
            .O(N__35492),
            .I(N__35396));
    Span4Mux_h I__7211 (
            .O(N__35489),
            .I(N__35393));
    Span4Mux_v I__7210 (
            .O(N__35484),
            .I(N__35386));
    Span4Mux_v I__7209 (
            .O(N__35481),
            .I(N__35386));
    Span4Mux_v I__7208 (
            .O(N__35472),
            .I(N__35386));
    InMux I__7207 (
            .O(N__35471),
            .I(N__35379));
    InMux I__7206 (
            .O(N__35468),
            .I(N__35379));
    InMux I__7205 (
            .O(N__35467),
            .I(N__35379));
    LocalMux I__7204 (
            .O(N__35452),
            .I(N__35372));
    LocalMux I__7203 (
            .O(N__35435),
            .I(N__35372));
    LocalMux I__7202 (
            .O(N__35430),
            .I(N__35372));
    InMux I__7201 (
            .O(N__35427),
            .I(N__35355));
    InMux I__7200 (
            .O(N__35426),
            .I(N__35355));
    InMux I__7199 (
            .O(N__35423),
            .I(N__35355));
    InMux I__7198 (
            .O(N__35422),
            .I(N__35355));
    InMux I__7197 (
            .O(N__35419),
            .I(N__35355));
    InMux I__7196 (
            .O(N__35418),
            .I(N__35355));
    InMux I__7195 (
            .O(N__35415),
            .I(N__35355));
    InMux I__7194 (
            .O(N__35414),
            .I(N__35355));
    InMux I__7193 (
            .O(N__35413),
            .I(N__35340));
    InMux I__7192 (
            .O(N__35410),
            .I(N__35340));
    InMux I__7191 (
            .O(N__35409),
            .I(N__35340));
    InMux I__7190 (
            .O(N__35406),
            .I(N__35340));
    InMux I__7189 (
            .O(N__35405),
            .I(N__35340));
    InMux I__7188 (
            .O(N__35402),
            .I(N__35340));
    InMux I__7187 (
            .O(N__35401),
            .I(N__35340));
    Span12Mux_s11_h I__7186 (
            .O(N__35396),
            .I(N__35337));
    Span4Mux_h I__7185 (
            .O(N__35393),
            .I(N__35334));
    Span4Mux_h I__7184 (
            .O(N__35386),
            .I(N__35331));
    LocalMux I__7183 (
            .O(N__35379),
            .I(N__35328));
    Span4Mux_v I__7182 (
            .O(N__35372),
            .I(N__35321));
    LocalMux I__7181 (
            .O(N__35355),
            .I(N__35321));
    LocalMux I__7180 (
            .O(N__35340),
            .I(N__35321));
    Span12Mux_v I__7179 (
            .O(N__35337),
            .I(N__35318));
    Span4Mux_h I__7178 (
            .O(N__35334),
            .I(N__35313));
    Span4Mux_h I__7177 (
            .O(N__35331),
            .I(N__35313));
    Span4Mux_v I__7176 (
            .O(N__35328),
            .I(N__35308));
    Span4Mux_v I__7175 (
            .O(N__35321),
            .I(N__35308));
    Odrv12 I__7174 (
            .O(N__35318),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7173 (
            .O(N__35313),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7172 (
            .O(N__35308),
            .I(CONSTANT_ONE_NET));
    InMux I__7171 (
            .O(N__35301),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__7170 (
            .O(N__35298),
            .I(N__35291));
    InMux I__7169 (
            .O(N__35297),
            .I(N__35291));
    CascadeMux I__7168 (
            .O(N__35296),
            .I(N__35279));
    LocalMux I__7167 (
            .O(N__35291),
            .I(N__35273));
    InMux I__7166 (
            .O(N__35290),
            .I(N__35258));
    InMux I__7165 (
            .O(N__35289),
            .I(N__35258));
    InMux I__7164 (
            .O(N__35288),
            .I(N__35258));
    InMux I__7163 (
            .O(N__35287),
            .I(N__35258));
    InMux I__7162 (
            .O(N__35286),
            .I(N__35258));
    InMux I__7161 (
            .O(N__35285),
            .I(N__35258));
    InMux I__7160 (
            .O(N__35284),
            .I(N__35258));
    InMux I__7159 (
            .O(N__35283),
            .I(N__35253));
    InMux I__7158 (
            .O(N__35282),
            .I(N__35253));
    InMux I__7157 (
            .O(N__35279),
            .I(N__35250));
    InMux I__7156 (
            .O(N__35278),
            .I(N__35243));
    InMux I__7155 (
            .O(N__35277),
            .I(N__35243));
    InMux I__7154 (
            .O(N__35276),
            .I(N__35243));
    Span4Mux_h I__7153 (
            .O(N__35273),
            .I(N__35238));
    LocalMux I__7152 (
            .O(N__35258),
            .I(N__35238));
    LocalMux I__7151 (
            .O(N__35253),
            .I(N__35235));
    LocalMux I__7150 (
            .O(N__35250),
            .I(N__35230));
    LocalMux I__7149 (
            .O(N__35243),
            .I(N__35230));
    Span4Mux_h I__7148 (
            .O(N__35238),
            .I(N__35227));
    Span4Mux_h I__7147 (
            .O(N__35235),
            .I(N__35224));
    Span4Mux_h I__7146 (
            .O(N__35230),
            .I(N__35219));
    Span4Mux_v I__7145 (
            .O(N__35227),
            .I(N__35219));
    Odrv4 I__7144 (
            .O(N__35224),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__7143 (
            .O(N__35219),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__7142 (
            .O(N__35214),
            .I(N__35211));
    LocalMux I__7141 (
            .O(N__35211),
            .I(N__35205));
    InMux I__7140 (
            .O(N__35210),
            .I(N__35202));
    InMux I__7139 (
            .O(N__35209),
            .I(N__35197));
    InMux I__7138 (
            .O(N__35208),
            .I(N__35197));
    Span12Mux_v I__7137 (
            .O(N__35205),
            .I(N__35194));
    LocalMux I__7136 (
            .O(N__35202),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__7135 (
            .O(N__35197),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv12 I__7134 (
            .O(N__35194),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__7133 (
            .O(N__35187),
            .I(N__35183));
    InMux I__7132 (
            .O(N__35186),
            .I(N__35179));
    LocalMux I__7131 (
            .O(N__35183),
            .I(N__35176));
    InMux I__7130 (
            .O(N__35182),
            .I(N__35173));
    LocalMux I__7129 (
            .O(N__35179),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__7128 (
            .O(N__35176),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__7127 (
            .O(N__35173),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__7126 (
            .O(N__35166),
            .I(N__35162));
    InMux I__7125 (
            .O(N__35165),
            .I(N__35158));
    LocalMux I__7124 (
            .O(N__35162),
            .I(N__35155));
    InMux I__7123 (
            .O(N__35161),
            .I(N__35152));
    LocalMux I__7122 (
            .O(N__35158),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__7121 (
            .O(N__35155),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__7120 (
            .O(N__35152),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__7119 (
            .O(N__35145),
            .I(N__35140));
    InMux I__7118 (
            .O(N__35144),
            .I(N__35137));
    InMux I__7117 (
            .O(N__35143),
            .I(N__35134));
    LocalMux I__7116 (
            .O(N__35140),
            .I(N__35131));
    LocalMux I__7115 (
            .O(N__35137),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__7114 (
            .O(N__35134),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__7113 (
            .O(N__35131),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__7112 (
            .O(N__35124),
            .I(N__35120));
    InMux I__7111 (
            .O(N__35123),
            .I(N__35116));
    LocalMux I__7110 (
            .O(N__35120),
            .I(N__35113));
    InMux I__7109 (
            .O(N__35119),
            .I(N__35110));
    LocalMux I__7108 (
            .O(N__35116),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__7107 (
            .O(N__35113),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__7106 (
            .O(N__35110),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__7105 (
            .O(N__35103),
            .I(N__35099));
    InMux I__7104 (
            .O(N__35102),
            .I(N__35095));
    LocalMux I__7103 (
            .O(N__35099),
            .I(N__35092));
    InMux I__7102 (
            .O(N__35098),
            .I(N__35089));
    LocalMux I__7101 (
            .O(N__35095),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__7100 (
            .O(N__35092),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__7099 (
            .O(N__35089),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__7098 (
            .O(N__35082),
            .I(N__35077));
    InMux I__7097 (
            .O(N__35081),
            .I(N__35074));
    InMux I__7096 (
            .O(N__35080),
            .I(N__35071));
    LocalMux I__7095 (
            .O(N__35077),
            .I(N__35068));
    LocalMux I__7094 (
            .O(N__35074),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__7093 (
            .O(N__35071),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__7092 (
            .O(N__35068),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__7091 (
            .O(N__35061),
            .I(N__35056));
    InMux I__7090 (
            .O(N__35060),
            .I(N__35053));
    InMux I__7089 (
            .O(N__35059),
            .I(N__35050));
    LocalMux I__7088 (
            .O(N__35056),
            .I(N__35047));
    LocalMux I__7087 (
            .O(N__35053),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__7086 (
            .O(N__35050),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__7085 (
            .O(N__35047),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    CascadeMux I__7084 (
            .O(N__35040),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__7083 (
            .O(N__35037),
            .I(N__35032));
    InMux I__7082 (
            .O(N__35036),
            .I(N__35029));
    InMux I__7081 (
            .O(N__35035),
            .I(N__35026));
    LocalMux I__7080 (
            .O(N__35032),
            .I(N__35023));
    LocalMux I__7079 (
            .O(N__35029),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__7078 (
            .O(N__35026),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__7077 (
            .O(N__35023),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__7076 (
            .O(N__35016),
            .I(N__35013));
    LocalMux I__7075 (
            .O(N__35013),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    InMux I__7074 (
            .O(N__35010),
            .I(N__35005));
    InMux I__7073 (
            .O(N__35009),
            .I(N__35002));
    InMux I__7072 (
            .O(N__35008),
            .I(N__34999));
    LocalMux I__7071 (
            .O(N__35005),
            .I(N__34996));
    LocalMux I__7070 (
            .O(N__35002),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__7069 (
            .O(N__34999),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__7068 (
            .O(N__34996),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    CascadeMux I__7067 (
            .O(N__34989),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__7066 (
            .O(N__34986),
            .I(N__34981));
    InMux I__7065 (
            .O(N__34985),
            .I(N__34978));
    InMux I__7064 (
            .O(N__34984),
            .I(N__34975));
    LocalMux I__7063 (
            .O(N__34981),
            .I(N__34972));
    LocalMux I__7062 (
            .O(N__34978),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__7061 (
            .O(N__34975),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv12 I__7060 (
            .O(N__34972),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__7059 (
            .O(N__34965),
            .I(N__34947));
    InMux I__7058 (
            .O(N__34964),
            .I(N__34947));
    InMux I__7057 (
            .O(N__34963),
            .I(N__34947));
    InMux I__7056 (
            .O(N__34962),
            .I(N__34947));
    InMux I__7055 (
            .O(N__34961),
            .I(N__34942));
    InMux I__7054 (
            .O(N__34960),
            .I(N__34942));
    InMux I__7053 (
            .O(N__34959),
            .I(N__34933));
    InMux I__7052 (
            .O(N__34958),
            .I(N__34933));
    InMux I__7051 (
            .O(N__34957),
            .I(N__34933));
    InMux I__7050 (
            .O(N__34956),
            .I(N__34933));
    LocalMux I__7049 (
            .O(N__34947),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__7048 (
            .O(N__34942),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__7047 (
            .O(N__34933),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__7046 (
            .O(N__34926),
            .I(N__34923));
    LocalMux I__7045 (
            .O(N__34923),
            .I(N__34920));
    Odrv4 I__7044 (
            .O(N__34920),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__7043 (
            .O(N__34917),
            .I(N__34914));
    LocalMux I__7042 (
            .O(N__34914),
            .I(N__34911));
    Odrv4 I__7041 (
            .O(N__34911),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    CascadeMux I__7040 (
            .O(N__34908),
            .I(N__34905));
    InMux I__7039 (
            .O(N__34905),
            .I(N__34902));
    LocalMux I__7038 (
            .O(N__34902),
            .I(N__34899));
    Odrv4 I__7037 (
            .O(N__34899),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__7036 (
            .O(N__34896),
            .I(N__34893));
    InMux I__7035 (
            .O(N__34893),
            .I(N__34890));
    LocalMux I__7034 (
            .O(N__34890),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__7033 (
            .O(N__34887),
            .I(N__34884));
    LocalMux I__7032 (
            .O(N__34884),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    InMux I__7031 (
            .O(N__34881),
            .I(N__34878));
    LocalMux I__7030 (
            .O(N__34878),
            .I(N__34875));
    Odrv4 I__7029 (
            .O(N__34875),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__7028 (
            .O(N__34872),
            .I(N__34869));
    InMux I__7027 (
            .O(N__34869),
            .I(N__34866));
    LocalMux I__7026 (
            .O(N__34866),
            .I(N__34863));
    Odrv4 I__7025 (
            .O(N__34863),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__7024 (
            .O(N__34860),
            .I(N__34857));
    InMux I__7023 (
            .O(N__34857),
            .I(N__34854));
    LocalMux I__7022 (
            .O(N__34854),
            .I(N__34851));
    Odrv4 I__7021 (
            .O(N__34851),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__7020 (
            .O(N__34848),
            .I(N__34845));
    LocalMux I__7019 (
            .O(N__34845),
            .I(N__34842));
    Odrv12 I__7018 (
            .O(N__34842),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__7017 (
            .O(N__34839),
            .I(N__34836));
    LocalMux I__7016 (
            .O(N__34836),
            .I(N__34833));
    Span4Mux_h I__7015 (
            .O(N__34833),
            .I(N__34830));
    Odrv4 I__7014 (
            .O(N__34830),
            .I(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ));
    InMux I__7013 (
            .O(N__34827),
            .I(N__34824));
    LocalMux I__7012 (
            .O(N__34824),
            .I(N__34821));
    Span4Mux_h I__7011 (
            .O(N__34821),
            .I(N__34818));
    Odrv4 I__7010 (
            .O(N__34818),
            .I(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ));
    InMux I__7009 (
            .O(N__34815),
            .I(N__34812));
    LocalMux I__7008 (
            .O(N__34812),
            .I(N__34809));
    Span4Mux_v I__7007 (
            .O(N__34809),
            .I(N__34806));
    Odrv4 I__7006 (
            .O(N__34806),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__7005 (
            .O(N__34803),
            .I(N__34800));
    LocalMux I__7004 (
            .O(N__34800),
            .I(N__34797));
    Span4Mux_v I__7003 (
            .O(N__34797),
            .I(N__34794));
    Odrv4 I__7002 (
            .O(N__34794),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    CascadeMux I__7001 (
            .O(N__34791),
            .I(N__34788));
    InMux I__7000 (
            .O(N__34788),
            .I(N__34785));
    LocalMux I__6999 (
            .O(N__34785),
            .I(N__34782));
    Span4Mux_h I__6998 (
            .O(N__34782),
            .I(N__34779));
    Odrv4 I__6997 (
            .O(N__34779),
            .I(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ));
    CascadeMux I__6996 (
            .O(N__34776),
            .I(N__34773));
    InMux I__6995 (
            .O(N__34773),
            .I(N__34770));
    LocalMux I__6994 (
            .O(N__34770),
            .I(N__34767));
    Span4Mux_v I__6993 (
            .O(N__34767),
            .I(N__34764));
    Odrv4 I__6992 (
            .O(N__34764),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    CascadeMux I__6991 (
            .O(N__34761),
            .I(N__34758));
    InMux I__6990 (
            .O(N__34758),
            .I(N__34754));
    InMux I__6989 (
            .O(N__34757),
            .I(N__34751));
    LocalMux I__6988 (
            .O(N__34754),
            .I(N__34748));
    LocalMux I__6987 (
            .O(N__34751),
            .I(N__34745));
    Span4Mux_v I__6986 (
            .O(N__34748),
            .I(N__34742));
    Odrv12 I__6985 (
            .O(N__34745),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv4 I__6984 (
            .O(N__34742),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__6983 (
            .O(N__34737),
            .I(N__34734));
    LocalMux I__6982 (
            .O(N__34734),
            .I(N__34731));
    Odrv12 I__6981 (
            .O(N__34731),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__6980 (
            .O(N__34728),
            .I(N__34725));
    InMux I__6979 (
            .O(N__34725),
            .I(N__34722));
    LocalMux I__6978 (
            .O(N__34722),
            .I(N__34719));
    Span4Mux_v I__6977 (
            .O(N__34719),
            .I(N__34716));
    Odrv4 I__6976 (
            .O(N__34716),
            .I(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ));
    CascadeMux I__6975 (
            .O(N__34713),
            .I(N__34710));
    InMux I__6974 (
            .O(N__34710),
            .I(N__34707));
    LocalMux I__6973 (
            .O(N__34707),
            .I(N__34704));
    Span4Mux_v I__6972 (
            .O(N__34704),
            .I(N__34701));
    Odrv4 I__6971 (
            .O(N__34701),
            .I(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ));
    InMux I__6970 (
            .O(N__34698),
            .I(N__34695));
    LocalMux I__6969 (
            .O(N__34695),
            .I(N__34692));
    Span4Mux_v I__6968 (
            .O(N__34692),
            .I(N__34689));
    Odrv4 I__6967 (
            .O(N__34689),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    CascadeMux I__6966 (
            .O(N__34686),
            .I(N__34683));
    InMux I__6965 (
            .O(N__34683),
            .I(N__34680));
    LocalMux I__6964 (
            .O(N__34680),
            .I(N__34677));
    Span4Mux_v I__6963 (
            .O(N__34677),
            .I(N__34674));
    Odrv4 I__6962 (
            .O(N__34674),
            .I(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ));
    InMux I__6961 (
            .O(N__34671),
            .I(N__34668));
    LocalMux I__6960 (
            .O(N__34668),
            .I(N__34665));
    Span4Mux_v I__6959 (
            .O(N__34665),
            .I(N__34662));
    Odrv4 I__6958 (
            .O(N__34662),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    CascadeMux I__6957 (
            .O(N__34659),
            .I(N__34656));
    InMux I__6956 (
            .O(N__34656),
            .I(N__34653));
    LocalMux I__6955 (
            .O(N__34653),
            .I(N__34650));
    Span4Mux_v I__6954 (
            .O(N__34650),
            .I(N__34647));
    Odrv4 I__6953 (
            .O(N__34647),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__6952 (
            .O(N__34644),
            .I(N__34641));
    LocalMux I__6951 (
            .O(N__34641),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ));
    InMux I__6950 (
            .O(N__34638),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ));
    InMux I__6949 (
            .O(N__34635),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    CascadeMux I__6948 (
            .O(N__34632),
            .I(N__34629));
    InMux I__6947 (
            .O(N__34629),
            .I(N__34626));
    LocalMux I__6946 (
            .O(N__34626),
            .I(N__34623));
    Span4Mux_v I__6945 (
            .O(N__34623),
            .I(N__34620));
    Odrv4 I__6944 (
            .O(N__34620),
            .I(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ));
    CascadeMux I__6943 (
            .O(N__34617),
            .I(N__34614));
    InMux I__6942 (
            .O(N__34614),
            .I(N__34611));
    LocalMux I__6941 (
            .O(N__34611),
            .I(N__34608));
    Span4Mux_v I__6940 (
            .O(N__34608),
            .I(N__34605));
    Odrv4 I__6939 (
            .O(N__34605),
            .I(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ));
    CascadeMux I__6938 (
            .O(N__34602),
            .I(N__34599));
    InMux I__6937 (
            .O(N__34599),
            .I(N__34596));
    LocalMux I__6936 (
            .O(N__34596),
            .I(N__34593));
    Span4Mux_v I__6935 (
            .O(N__34593),
            .I(N__34590));
    Odrv4 I__6934 (
            .O(N__34590),
            .I(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ));
    CascadeMux I__6933 (
            .O(N__34587),
            .I(N__34584));
    InMux I__6932 (
            .O(N__34584),
            .I(N__34581));
    LocalMux I__6931 (
            .O(N__34581),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__6930 (
            .O(N__34578),
            .I(N__34575));
    InMux I__6929 (
            .O(N__34575),
            .I(N__34572));
    LocalMux I__6928 (
            .O(N__34572),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__6927 (
            .O(N__34569),
            .I(N__34566));
    LocalMux I__6926 (
            .O(N__34566),
            .I(N__34563));
    Odrv4 I__6925 (
            .O(N__34563),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ));
    CascadeMux I__6924 (
            .O(N__34560),
            .I(N__34557));
    InMux I__6923 (
            .O(N__34557),
            .I(N__34554));
    LocalMux I__6922 (
            .O(N__34554),
            .I(N__34551));
    Odrv4 I__6921 (
            .O(N__34551),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt22 ));
    CascadeMux I__6920 (
            .O(N__34548),
            .I(N__34545));
    InMux I__6919 (
            .O(N__34545),
            .I(N__34542));
    LocalMux I__6918 (
            .O(N__34542),
            .I(N__34539));
    Odrv4 I__6917 (
            .O(N__34539),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__6916 (
            .O(N__34536),
            .I(N__34533));
    LocalMux I__6915 (
            .O(N__34533),
            .I(N__34530));
    Odrv4 I__6914 (
            .O(N__34530),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__6913 (
            .O(N__34527),
            .I(N__34524));
    InMux I__6912 (
            .O(N__34524),
            .I(N__34521));
    LocalMux I__6911 (
            .O(N__34521),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__6910 (
            .O(N__34518),
            .I(N__34515));
    LocalMux I__6909 (
            .O(N__34515),
            .I(N__34512));
    Span4Mux_h I__6908 (
            .O(N__34512),
            .I(N__34509));
    Odrv4 I__6907 (
            .O(N__34509),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__6906 (
            .O(N__34506),
            .I(N__34503));
    InMux I__6905 (
            .O(N__34503),
            .I(N__34500));
    LocalMux I__6904 (
            .O(N__34500),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__6903 (
            .O(N__34497),
            .I(N__34494));
    LocalMux I__6902 (
            .O(N__34494),
            .I(N__34491));
    Odrv12 I__6901 (
            .O(N__34491),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__6900 (
            .O(N__34488),
            .I(N__34485));
    InMux I__6899 (
            .O(N__34485),
            .I(N__34482));
    LocalMux I__6898 (
            .O(N__34482),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__6897 (
            .O(N__34479),
            .I(N__34476));
    InMux I__6896 (
            .O(N__34476),
            .I(N__34473));
    LocalMux I__6895 (
            .O(N__34473),
            .I(N__34470));
    Odrv4 I__6894 (
            .O(N__34470),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    InMux I__6893 (
            .O(N__34467),
            .I(N__34464));
    LocalMux I__6892 (
            .O(N__34464),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__6891 (
            .O(N__34461),
            .I(N__34458));
    LocalMux I__6890 (
            .O(N__34458),
            .I(N__34455));
    Odrv4 I__6889 (
            .O(N__34455),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__6888 (
            .O(N__34452),
            .I(N__34449));
    InMux I__6887 (
            .O(N__34449),
            .I(N__34446));
    LocalMux I__6886 (
            .O(N__34446),
            .I(N__34443));
    Odrv4 I__6885 (
            .O(N__34443),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__6884 (
            .O(N__34440),
            .I(N__34437));
    LocalMux I__6883 (
            .O(N__34437),
            .I(N__34434));
    Odrv4 I__6882 (
            .O(N__34434),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__6881 (
            .O(N__34431),
            .I(N__34428));
    InMux I__6880 (
            .O(N__34428),
            .I(N__34425));
    LocalMux I__6879 (
            .O(N__34425),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__6878 (
            .O(N__34422),
            .I(N__34419));
    InMux I__6877 (
            .O(N__34419),
            .I(N__34416));
    LocalMux I__6876 (
            .O(N__34416),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__6875 (
            .O(N__34413),
            .I(N__34410));
    LocalMux I__6874 (
            .O(N__34410),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__6873 (
            .O(N__34407),
            .I(N__34404));
    LocalMux I__6872 (
            .O(N__34404),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    InMux I__6871 (
            .O(N__34401),
            .I(N__34398));
    LocalMux I__6870 (
            .O(N__34398),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ));
    CascadeMux I__6869 (
            .O(N__34395),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21_cascade_));
    CascadeMux I__6868 (
            .O(N__34392),
            .I(N__34389));
    InMux I__6867 (
            .O(N__34389),
            .I(N__34386));
    LocalMux I__6866 (
            .O(N__34386),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__6865 (
            .O(N__34383),
            .I(N__34380));
    LocalMux I__6864 (
            .O(N__34380),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__6863 (
            .O(N__34377),
            .I(N__34374));
    InMux I__6862 (
            .O(N__34374),
            .I(N__34371));
    LocalMux I__6861 (
            .O(N__34371),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__6860 (
            .O(N__34368),
            .I(N__34365));
    InMux I__6859 (
            .O(N__34365),
            .I(N__34362));
    LocalMux I__6858 (
            .O(N__34362),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__6857 (
            .O(N__34359),
            .I(N__34356));
    InMux I__6856 (
            .O(N__34356),
            .I(N__34353));
    LocalMux I__6855 (
            .O(N__34353),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__6854 (
            .O(N__34350),
            .I(N__34322));
    InMux I__6853 (
            .O(N__34349),
            .I(N__34322));
    InMux I__6852 (
            .O(N__34348),
            .I(N__34322));
    InMux I__6851 (
            .O(N__34347),
            .I(N__34322));
    InMux I__6850 (
            .O(N__34346),
            .I(N__34313));
    InMux I__6849 (
            .O(N__34345),
            .I(N__34313));
    InMux I__6848 (
            .O(N__34344),
            .I(N__34313));
    InMux I__6847 (
            .O(N__34343),
            .I(N__34313));
    InMux I__6846 (
            .O(N__34342),
            .I(N__34294));
    InMux I__6845 (
            .O(N__34341),
            .I(N__34294));
    InMux I__6844 (
            .O(N__34340),
            .I(N__34294));
    InMux I__6843 (
            .O(N__34339),
            .I(N__34294));
    InMux I__6842 (
            .O(N__34338),
            .I(N__34285));
    InMux I__6841 (
            .O(N__34337),
            .I(N__34285));
    InMux I__6840 (
            .O(N__34336),
            .I(N__34285));
    InMux I__6839 (
            .O(N__34335),
            .I(N__34285));
    InMux I__6838 (
            .O(N__34334),
            .I(N__34276));
    InMux I__6837 (
            .O(N__34333),
            .I(N__34276));
    InMux I__6836 (
            .O(N__34332),
            .I(N__34276));
    InMux I__6835 (
            .O(N__34331),
            .I(N__34276));
    LocalMux I__6834 (
            .O(N__34322),
            .I(N__34271));
    LocalMux I__6833 (
            .O(N__34313),
            .I(N__34271));
    InMux I__6832 (
            .O(N__34312),
            .I(N__34266));
    InMux I__6831 (
            .O(N__34311),
            .I(N__34266));
    InMux I__6830 (
            .O(N__34310),
            .I(N__34257));
    InMux I__6829 (
            .O(N__34309),
            .I(N__34257));
    InMux I__6828 (
            .O(N__34308),
            .I(N__34257));
    InMux I__6827 (
            .O(N__34307),
            .I(N__34257));
    InMux I__6826 (
            .O(N__34306),
            .I(N__34248));
    InMux I__6825 (
            .O(N__34305),
            .I(N__34248));
    InMux I__6824 (
            .O(N__34304),
            .I(N__34248));
    InMux I__6823 (
            .O(N__34303),
            .I(N__34248));
    LocalMux I__6822 (
            .O(N__34294),
            .I(N__34245));
    LocalMux I__6821 (
            .O(N__34285),
            .I(N__34238));
    LocalMux I__6820 (
            .O(N__34276),
            .I(N__34238));
    Span4Mux_h I__6819 (
            .O(N__34271),
            .I(N__34238));
    LocalMux I__6818 (
            .O(N__34266),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__6817 (
            .O(N__34257),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__6816 (
            .O(N__34248),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv12 I__6815 (
            .O(N__34245),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__6814 (
            .O(N__34238),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    CascadeMux I__6813 (
            .O(N__34227),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_ ));
    InMux I__6812 (
            .O(N__34224),
            .I(N__34221));
    LocalMux I__6811 (
            .O(N__34221),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ));
    CascadeMux I__6810 (
            .O(N__34218),
            .I(N__34214));
    CascadeMux I__6809 (
            .O(N__34217),
            .I(N__34211));
    InMux I__6808 (
            .O(N__34214),
            .I(N__34205));
    InMux I__6807 (
            .O(N__34211),
            .I(N__34205));
    InMux I__6806 (
            .O(N__34210),
            .I(N__34202));
    LocalMux I__6805 (
            .O(N__34205),
            .I(N__34199));
    LocalMux I__6804 (
            .O(N__34202),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv4 I__6803 (
            .O(N__34199),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__6802 (
            .O(N__34194),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__6801 (
            .O(N__34191),
            .I(N__34184));
    InMux I__6800 (
            .O(N__34190),
            .I(N__34184));
    InMux I__6799 (
            .O(N__34189),
            .I(N__34181));
    LocalMux I__6798 (
            .O(N__34184),
            .I(N__34178));
    LocalMux I__6797 (
            .O(N__34181),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__6796 (
            .O(N__34178),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__6795 (
            .O(N__34173),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    CascadeMux I__6794 (
            .O(N__34170),
            .I(N__34166));
    InMux I__6793 (
            .O(N__34169),
            .I(N__34163));
    InMux I__6792 (
            .O(N__34166),
            .I(N__34159));
    LocalMux I__6791 (
            .O(N__34163),
            .I(N__34156));
    InMux I__6790 (
            .O(N__34162),
            .I(N__34153));
    LocalMux I__6789 (
            .O(N__34159),
            .I(N__34148));
    Span4Mux_h I__6788 (
            .O(N__34156),
            .I(N__34148));
    LocalMux I__6787 (
            .O(N__34153),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__6786 (
            .O(N__34148),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__6785 (
            .O(N__34143),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__6784 (
            .O(N__34140),
            .I(N__34136));
    CascadeMux I__6783 (
            .O(N__34139),
            .I(N__34132));
    LocalMux I__6782 (
            .O(N__34136),
            .I(N__34129));
    InMux I__6781 (
            .O(N__34135),
            .I(N__34126));
    InMux I__6780 (
            .O(N__34132),
            .I(N__34123));
    Span4Mux_v I__6779 (
            .O(N__34129),
            .I(N__34120));
    LocalMux I__6778 (
            .O(N__34126),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__6777 (
            .O(N__34123),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__6776 (
            .O(N__34120),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__6775 (
            .O(N__34113),
            .I(bfn_14_8_0_));
    CascadeMux I__6774 (
            .O(N__34110),
            .I(N__34107));
    InMux I__6773 (
            .O(N__34107),
            .I(N__34104));
    LocalMux I__6772 (
            .O(N__34104),
            .I(N__34100));
    InMux I__6771 (
            .O(N__34103),
            .I(N__34096));
    Span4Mux_h I__6770 (
            .O(N__34100),
            .I(N__34093));
    InMux I__6769 (
            .O(N__34099),
            .I(N__34090));
    LocalMux I__6768 (
            .O(N__34096),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__6767 (
            .O(N__34093),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__6766 (
            .O(N__34090),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__6765 (
            .O(N__34083),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    CascadeMux I__6764 (
            .O(N__34080),
            .I(N__34076));
    CascadeMux I__6763 (
            .O(N__34079),
            .I(N__34073));
    InMux I__6762 (
            .O(N__34076),
            .I(N__34067));
    InMux I__6761 (
            .O(N__34073),
            .I(N__34067));
    InMux I__6760 (
            .O(N__34072),
            .I(N__34064));
    LocalMux I__6759 (
            .O(N__34067),
            .I(N__34061));
    LocalMux I__6758 (
            .O(N__34064),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv4 I__6757 (
            .O(N__34061),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__6756 (
            .O(N__34056),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__6755 (
            .O(N__34053),
            .I(N__34046));
    InMux I__6754 (
            .O(N__34052),
            .I(N__34046));
    InMux I__6753 (
            .O(N__34051),
            .I(N__34043));
    LocalMux I__6752 (
            .O(N__34046),
            .I(N__34040));
    LocalMux I__6751 (
            .O(N__34043),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__6750 (
            .O(N__34040),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__6749 (
            .O(N__34035),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__6748 (
            .O(N__34032),
            .I(N__34028));
    InMux I__6747 (
            .O(N__34031),
            .I(N__34025));
    LocalMux I__6746 (
            .O(N__34028),
            .I(N__34022));
    LocalMux I__6745 (
            .O(N__34025),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv4 I__6744 (
            .O(N__34022),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__6743 (
            .O(N__34017),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__6742 (
            .O(N__34014),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CascadeMux I__6741 (
            .O(N__34011),
            .I(N__34008));
    InMux I__6740 (
            .O(N__34008),
            .I(N__34004));
    InMux I__6739 (
            .O(N__34007),
            .I(N__34001));
    LocalMux I__6738 (
            .O(N__34004),
            .I(N__33998));
    LocalMux I__6737 (
            .O(N__34001),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__6736 (
            .O(N__33998),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__6735 (
            .O(N__33993),
            .I(N__33988));
    CEMux I__6734 (
            .O(N__33992),
            .I(N__33985));
    CEMux I__6733 (
            .O(N__33991),
            .I(N__33981));
    LocalMux I__6732 (
            .O(N__33988),
            .I(N__33978));
    LocalMux I__6731 (
            .O(N__33985),
            .I(N__33975));
    CEMux I__6730 (
            .O(N__33984),
            .I(N__33972));
    LocalMux I__6729 (
            .O(N__33981),
            .I(N__33969));
    Span4Mux_v I__6728 (
            .O(N__33978),
            .I(N__33962));
    Span4Mux_v I__6727 (
            .O(N__33975),
            .I(N__33962));
    LocalMux I__6726 (
            .O(N__33972),
            .I(N__33962));
    Span4Mux_v I__6725 (
            .O(N__33969),
            .I(N__33959));
    Span4Mux_v I__6724 (
            .O(N__33962),
            .I(N__33956));
    Span4Mux_v I__6723 (
            .O(N__33959),
            .I(N__33953));
    Span4Mux_v I__6722 (
            .O(N__33956),
            .I(N__33950));
    Span4Mux_v I__6721 (
            .O(N__33953),
            .I(N__33947));
    Span4Mux_v I__6720 (
            .O(N__33950),
            .I(N__33944));
    Odrv4 I__6719 (
            .O(N__33947),
            .I(\delay_measurement_inst.delay_tr_timer.N_201_i ));
    Odrv4 I__6718 (
            .O(N__33944),
            .I(\delay_measurement_inst.delay_tr_timer.N_201_i ));
    CascadeMux I__6717 (
            .O(N__33939),
            .I(N__33935));
    CascadeMux I__6716 (
            .O(N__33938),
            .I(N__33932));
    InMux I__6715 (
            .O(N__33935),
            .I(N__33926));
    InMux I__6714 (
            .O(N__33932),
            .I(N__33926));
    InMux I__6713 (
            .O(N__33931),
            .I(N__33923));
    LocalMux I__6712 (
            .O(N__33926),
            .I(N__33920));
    LocalMux I__6711 (
            .O(N__33923),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv4 I__6710 (
            .O(N__33920),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__6709 (
            .O(N__33915),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    CascadeMux I__6708 (
            .O(N__33912),
            .I(N__33908));
    CascadeMux I__6707 (
            .O(N__33911),
            .I(N__33905));
    InMux I__6706 (
            .O(N__33908),
            .I(N__33900));
    InMux I__6705 (
            .O(N__33905),
            .I(N__33900));
    LocalMux I__6704 (
            .O(N__33900),
            .I(N__33896));
    InMux I__6703 (
            .O(N__33899),
            .I(N__33893));
    Span4Mux_h I__6702 (
            .O(N__33896),
            .I(N__33890));
    LocalMux I__6701 (
            .O(N__33893),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__6700 (
            .O(N__33890),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__6699 (
            .O(N__33885),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__6698 (
            .O(N__33882),
            .I(N__33878));
    InMux I__6697 (
            .O(N__33881),
            .I(N__33875));
    InMux I__6696 (
            .O(N__33878),
            .I(N__33871));
    LocalMux I__6695 (
            .O(N__33875),
            .I(N__33868));
    InMux I__6694 (
            .O(N__33874),
            .I(N__33865));
    LocalMux I__6693 (
            .O(N__33871),
            .I(N__33860));
    Span4Mux_h I__6692 (
            .O(N__33868),
            .I(N__33860));
    LocalMux I__6691 (
            .O(N__33865),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__6690 (
            .O(N__33860),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__6689 (
            .O(N__33855),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    CascadeMux I__6688 (
            .O(N__33852),
            .I(N__33849));
    InMux I__6687 (
            .O(N__33849),
            .I(N__33846));
    LocalMux I__6686 (
            .O(N__33846),
            .I(N__33841));
    InMux I__6685 (
            .O(N__33845),
            .I(N__33838));
    InMux I__6684 (
            .O(N__33844),
            .I(N__33835));
    Odrv4 I__6683 (
            .O(N__33841),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__6682 (
            .O(N__33838),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__6681 (
            .O(N__33835),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__6680 (
            .O(N__33828),
            .I(bfn_14_7_0_));
    CascadeMux I__6679 (
            .O(N__33825),
            .I(N__33822));
    InMux I__6678 (
            .O(N__33822),
            .I(N__33819));
    LocalMux I__6677 (
            .O(N__33819),
            .I(N__33815));
    InMux I__6676 (
            .O(N__33818),
            .I(N__33811));
    Span4Mux_h I__6675 (
            .O(N__33815),
            .I(N__33808));
    InMux I__6674 (
            .O(N__33814),
            .I(N__33805));
    LocalMux I__6673 (
            .O(N__33811),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__6672 (
            .O(N__33808),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__6671 (
            .O(N__33805),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__6670 (
            .O(N__33798),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__6669 (
            .O(N__33795),
            .I(N__33788));
    InMux I__6668 (
            .O(N__33794),
            .I(N__33788));
    InMux I__6667 (
            .O(N__33793),
            .I(N__33785));
    LocalMux I__6666 (
            .O(N__33788),
            .I(N__33782));
    LocalMux I__6665 (
            .O(N__33785),
            .I(N__33777));
    Span4Mux_v I__6664 (
            .O(N__33782),
            .I(N__33777));
    Odrv4 I__6663 (
            .O(N__33777),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__6662 (
            .O(N__33774),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__6661 (
            .O(N__33771),
            .I(N__33764));
    InMux I__6660 (
            .O(N__33770),
            .I(N__33764));
    InMux I__6659 (
            .O(N__33769),
            .I(N__33761));
    LocalMux I__6658 (
            .O(N__33764),
            .I(N__33758));
    LocalMux I__6657 (
            .O(N__33761),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__6656 (
            .O(N__33758),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__6655 (
            .O(N__33753),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    CascadeMux I__6654 (
            .O(N__33750),
            .I(N__33746));
    CascadeMux I__6653 (
            .O(N__33749),
            .I(N__33743));
    InMux I__6652 (
            .O(N__33746),
            .I(N__33738));
    InMux I__6651 (
            .O(N__33743),
            .I(N__33738));
    LocalMux I__6650 (
            .O(N__33738),
            .I(N__33734));
    InMux I__6649 (
            .O(N__33737),
            .I(N__33731));
    Span4Mux_h I__6648 (
            .O(N__33734),
            .I(N__33728));
    LocalMux I__6647 (
            .O(N__33731),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__6646 (
            .O(N__33728),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__6645 (
            .O(N__33723),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    CascadeMux I__6644 (
            .O(N__33720),
            .I(N__33716));
    CascadeMux I__6643 (
            .O(N__33719),
            .I(N__33713));
    InMux I__6642 (
            .O(N__33716),
            .I(N__33707));
    InMux I__6641 (
            .O(N__33713),
            .I(N__33707));
    InMux I__6640 (
            .O(N__33712),
            .I(N__33704));
    LocalMux I__6639 (
            .O(N__33707),
            .I(N__33701));
    LocalMux I__6638 (
            .O(N__33704),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__6637 (
            .O(N__33701),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__6636 (
            .O(N__33696),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    CascadeMux I__6635 (
            .O(N__33693),
            .I(N__33689));
    CascadeMux I__6634 (
            .O(N__33692),
            .I(N__33686));
    InMux I__6633 (
            .O(N__33689),
            .I(N__33681));
    InMux I__6632 (
            .O(N__33686),
            .I(N__33681));
    LocalMux I__6631 (
            .O(N__33681),
            .I(N__33677));
    InMux I__6630 (
            .O(N__33680),
            .I(N__33674));
    Span4Mux_h I__6629 (
            .O(N__33677),
            .I(N__33671));
    LocalMux I__6628 (
            .O(N__33674),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__6627 (
            .O(N__33671),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__6626 (
            .O(N__33666),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__6625 (
            .O(N__33663),
            .I(N__33660));
    InMux I__6624 (
            .O(N__33660),
            .I(N__33656));
    InMux I__6623 (
            .O(N__33659),
            .I(N__33653));
    LocalMux I__6622 (
            .O(N__33656),
            .I(N__33647));
    LocalMux I__6621 (
            .O(N__33653),
            .I(N__33647));
    InMux I__6620 (
            .O(N__33652),
            .I(N__33644));
    Span4Mux_h I__6619 (
            .O(N__33647),
            .I(N__33641));
    LocalMux I__6618 (
            .O(N__33644),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__6617 (
            .O(N__33641),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__6616 (
            .O(N__33636),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__6615 (
            .O(N__33633),
            .I(N__33630));
    LocalMux I__6614 (
            .O(N__33630),
            .I(N__33627));
    Span4Mux_h I__6613 (
            .O(N__33627),
            .I(N__33622));
    InMux I__6612 (
            .O(N__33626),
            .I(N__33619));
    InMux I__6611 (
            .O(N__33625),
            .I(N__33616));
    Odrv4 I__6610 (
            .O(N__33622),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__6609 (
            .O(N__33619),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__6608 (
            .O(N__33616),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__6607 (
            .O(N__33609),
            .I(bfn_14_6_0_));
    CascadeMux I__6606 (
            .O(N__33606),
            .I(N__33603));
    InMux I__6605 (
            .O(N__33603),
            .I(N__33600));
    LocalMux I__6604 (
            .O(N__33600),
            .I(N__33596));
    InMux I__6603 (
            .O(N__33599),
            .I(N__33592));
    Span4Mux_h I__6602 (
            .O(N__33596),
            .I(N__33589));
    InMux I__6601 (
            .O(N__33595),
            .I(N__33586));
    LocalMux I__6600 (
            .O(N__33592),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__6599 (
            .O(N__33589),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__6598 (
            .O(N__33586),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__6597 (
            .O(N__33579),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__6596 (
            .O(N__33576),
            .I(N__33572));
    CascadeMux I__6595 (
            .O(N__33575),
            .I(N__33569));
    InMux I__6594 (
            .O(N__33572),
            .I(N__33563));
    InMux I__6593 (
            .O(N__33569),
            .I(N__33563));
    InMux I__6592 (
            .O(N__33568),
            .I(N__33560));
    LocalMux I__6591 (
            .O(N__33563),
            .I(N__33557));
    LocalMux I__6590 (
            .O(N__33560),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__6589 (
            .O(N__33557),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__6588 (
            .O(N__33552),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__6587 (
            .O(N__33549),
            .I(N__33542));
    InMux I__6586 (
            .O(N__33548),
            .I(N__33542));
    InMux I__6585 (
            .O(N__33547),
            .I(N__33539));
    LocalMux I__6584 (
            .O(N__33542),
            .I(N__33536));
    LocalMux I__6583 (
            .O(N__33539),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__6582 (
            .O(N__33536),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__6581 (
            .O(N__33531),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__6580 (
            .O(N__33528),
            .I(N__33521));
    InMux I__6579 (
            .O(N__33527),
            .I(N__33521));
    InMux I__6578 (
            .O(N__33526),
            .I(N__33518));
    LocalMux I__6577 (
            .O(N__33521),
            .I(N__33515));
    LocalMux I__6576 (
            .O(N__33518),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv4 I__6575 (
            .O(N__33515),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__6574 (
            .O(N__33510),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    CascadeMux I__6573 (
            .O(N__33507),
            .I(N__33504));
    InMux I__6572 (
            .O(N__33504),
            .I(N__33501));
    LocalMux I__6571 (
            .O(N__33501),
            .I(\pwm_generator_inst.threshold_9 ));
    InMux I__6570 (
            .O(N__33498),
            .I(N__33495));
    LocalMux I__6569 (
            .O(N__33495),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__6568 (
            .O(N__33492),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__6567 (
            .O(N__33489),
            .I(N__33486));
    LocalMux I__6566 (
            .O(N__33486),
            .I(N__33483));
    Span4Mux_s2_v I__6565 (
            .O(N__33483),
            .I(N__33480));
    Sp12to4 I__6564 (
            .O(N__33480),
            .I(N__33477));
    Span12Mux_h I__6563 (
            .O(N__33477),
            .I(N__33474));
    Span12Mux_v I__6562 (
            .O(N__33474),
            .I(N__33471));
    Odrv12 I__6561 (
            .O(N__33471),
            .I(pwm_output_c));
    CascadeMux I__6560 (
            .O(N__33468),
            .I(N__33465));
    InMux I__6559 (
            .O(N__33465),
            .I(N__33462));
    LocalMux I__6558 (
            .O(N__33462),
            .I(N__33458));
    InMux I__6557 (
            .O(N__33461),
            .I(N__33454));
    Span4Mux_h I__6556 (
            .O(N__33458),
            .I(N__33450));
    InMux I__6555 (
            .O(N__33457),
            .I(N__33447));
    LocalMux I__6554 (
            .O(N__33454),
            .I(N__33444));
    InMux I__6553 (
            .O(N__33453),
            .I(N__33441));
    Span4Mux_v I__6552 (
            .O(N__33450),
            .I(N__33438));
    LocalMux I__6551 (
            .O(N__33447),
            .I(N__33433));
    Span12Mux_v I__6550 (
            .O(N__33444),
            .I(N__33433));
    LocalMux I__6549 (
            .O(N__33441),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__6548 (
            .O(N__33438),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__6547 (
            .O(N__33433),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__6546 (
            .O(N__33426),
            .I(N__33423));
    LocalMux I__6545 (
            .O(N__33423),
            .I(N__33420));
    Odrv4 I__6544 (
            .O(N__33420),
            .I(s2_phy_c));
    InMux I__6543 (
            .O(N__33417),
            .I(bfn_14_5_0_));
    CascadeMux I__6542 (
            .O(N__33414),
            .I(N__33411));
    InMux I__6541 (
            .O(N__33411),
            .I(N__33408));
    LocalMux I__6540 (
            .O(N__33408),
            .I(N__33403));
    InMux I__6539 (
            .O(N__33407),
            .I(N__33400));
    InMux I__6538 (
            .O(N__33406),
            .I(N__33397));
    Span4Mux_h I__6537 (
            .O(N__33403),
            .I(N__33394));
    LocalMux I__6536 (
            .O(N__33400),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__6535 (
            .O(N__33397),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__6534 (
            .O(N__33394),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__6533 (
            .O(N__33387),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CascadeMux I__6532 (
            .O(N__33384),
            .I(N__33381));
    InMux I__6531 (
            .O(N__33381),
            .I(N__33376));
    InMux I__6530 (
            .O(N__33380),
            .I(N__33373));
    InMux I__6529 (
            .O(N__33379),
            .I(N__33370));
    LocalMux I__6528 (
            .O(N__33376),
            .I(N__33365));
    LocalMux I__6527 (
            .O(N__33373),
            .I(N__33365));
    LocalMux I__6526 (
            .O(N__33370),
            .I(N__33360));
    Span4Mux_v I__6525 (
            .O(N__33365),
            .I(N__33360));
    Odrv4 I__6524 (
            .O(N__33360),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__6523 (
            .O(N__33357),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__6522 (
            .O(N__33354),
            .I(N__33347));
    InMux I__6521 (
            .O(N__33353),
            .I(N__33347));
    InMux I__6520 (
            .O(N__33352),
            .I(N__33344));
    LocalMux I__6519 (
            .O(N__33347),
            .I(N__33341));
    LocalMux I__6518 (
            .O(N__33344),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__6517 (
            .O(N__33341),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__6516 (
            .O(N__33336),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__6515 (
            .O(N__33333),
            .I(N__33326));
    InMux I__6514 (
            .O(N__33332),
            .I(N__33326));
    InMux I__6513 (
            .O(N__33331),
            .I(N__33323));
    LocalMux I__6512 (
            .O(N__33326),
            .I(N__33320));
    LocalMux I__6511 (
            .O(N__33323),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv4 I__6510 (
            .O(N__33320),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__6509 (
            .O(N__33315),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__6508 (
            .O(N__33312),
            .I(N__33309));
    InMux I__6507 (
            .O(N__33309),
            .I(N__33306));
    LocalMux I__6506 (
            .O(N__33306),
            .I(\pwm_generator_inst.un14_counter_1 ));
    InMux I__6505 (
            .O(N__33303),
            .I(N__33300));
    LocalMux I__6504 (
            .O(N__33300),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__6503 (
            .O(N__33297),
            .I(N__33294));
    InMux I__6502 (
            .O(N__33294),
            .I(N__33291));
    LocalMux I__6501 (
            .O(N__33291),
            .I(N__33288));
    Odrv12 I__6500 (
            .O(N__33288),
            .I(\pwm_generator_inst.threshold_2 ));
    InMux I__6499 (
            .O(N__33285),
            .I(N__33282));
    LocalMux I__6498 (
            .O(N__33282),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__6497 (
            .O(N__33279),
            .I(N__33276));
    InMux I__6496 (
            .O(N__33276),
            .I(N__33273));
    LocalMux I__6495 (
            .O(N__33273),
            .I(N__33270));
    Odrv4 I__6494 (
            .O(N__33270),
            .I(\pwm_generator_inst.threshold_3 ));
    InMux I__6493 (
            .O(N__33267),
            .I(N__33264));
    LocalMux I__6492 (
            .O(N__33264),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__6491 (
            .O(N__33261),
            .I(N__33258));
    InMux I__6490 (
            .O(N__33258),
            .I(N__33255));
    LocalMux I__6489 (
            .O(N__33255),
            .I(N__33252));
    Odrv12 I__6488 (
            .O(N__33252),
            .I(\pwm_generator_inst.threshold_4 ));
    InMux I__6487 (
            .O(N__33249),
            .I(N__33246));
    LocalMux I__6486 (
            .O(N__33246),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__6485 (
            .O(N__33243),
            .I(N__33240));
    InMux I__6484 (
            .O(N__33240),
            .I(N__33237));
    LocalMux I__6483 (
            .O(N__33237),
            .I(\pwm_generator_inst.threshold_5 ));
    InMux I__6482 (
            .O(N__33234),
            .I(N__33231));
    LocalMux I__6481 (
            .O(N__33231),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__6480 (
            .O(N__33228),
            .I(N__33225));
    InMux I__6479 (
            .O(N__33225),
            .I(N__33222));
    LocalMux I__6478 (
            .O(N__33222),
            .I(\pwm_generator_inst.un14_counter_6 ));
    InMux I__6477 (
            .O(N__33219),
            .I(N__33216));
    LocalMux I__6476 (
            .O(N__33216),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__6475 (
            .O(N__33213),
            .I(N__33210));
    InMux I__6474 (
            .O(N__33210),
            .I(N__33207));
    LocalMux I__6473 (
            .O(N__33207),
            .I(\pwm_generator_inst.un14_counter_7 ));
    InMux I__6472 (
            .O(N__33204),
            .I(N__33201));
    LocalMux I__6471 (
            .O(N__33201),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__6470 (
            .O(N__33198),
            .I(N__33195));
    InMux I__6469 (
            .O(N__33195),
            .I(N__33192));
    LocalMux I__6468 (
            .O(N__33192),
            .I(N__33189));
    Odrv4 I__6467 (
            .O(N__33189),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__6466 (
            .O(N__33186),
            .I(N__33183));
    LocalMux I__6465 (
            .O(N__33183),
            .I(\pwm_generator_inst.counter_i_8 ));
    InMux I__6464 (
            .O(N__33180),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__6463 (
            .O(N__33177),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__6462 (
            .O(N__33174),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__6461 (
            .O(N__33171),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__6460 (
            .O(N__33168),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__6459 (
            .O(N__33165),
            .I(bfn_13_23_0_));
    InMux I__6458 (
            .O(N__33162),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__6457 (
            .O(N__33159),
            .I(N__33156));
    LocalMux I__6456 (
            .O(N__33156),
            .I(N__33152));
    InMux I__6455 (
            .O(N__33155),
            .I(N__33148));
    Span12Mux_v I__6454 (
            .O(N__33152),
            .I(N__33145));
    InMux I__6453 (
            .O(N__33151),
            .I(N__33142));
    LocalMux I__6452 (
            .O(N__33148),
            .I(N__33139));
    Odrv12 I__6451 (
            .O(N__33145),
            .I(il_min_comp1_D2));
    LocalMux I__6450 (
            .O(N__33142),
            .I(il_min_comp1_D2));
    Odrv12 I__6449 (
            .O(N__33139),
            .I(il_min_comp1_D2));
    InMux I__6448 (
            .O(N__33132),
            .I(N__33128));
    CascadeMux I__6447 (
            .O(N__33131),
            .I(N__33125));
    LocalMux I__6446 (
            .O(N__33128),
            .I(N__33122));
    InMux I__6445 (
            .O(N__33125),
            .I(N__33119));
    Span4Mux_v I__6444 (
            .O(N__33122),
            .I(N__33116));
    LocalMux I__6443 (
            .O(N__33119),
            .I(N__33113));
    Span4Mux_v I__6442 (
            .O(N__33116),
            .I(N__33110));
    Span12Mux_s7_v I__6441 (
            .O(N__33113),
            .I(N__33107));
    Odrv4 I__6440 (
            .O(N__33110),
            .I(\phase_controller_inst1.state_RNIE87FZ0Z_2 ));
    Odrv12 I__6439 (
            .O(N__33107),
            .I(\phase_controller_inst1.state_RNIE87FZ0Z_2 ));
    InMux I__6438 (
            .O(N__33102),
            .I(N__33099));
    LocalMux I__6437 (
            .O(N__33099),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__6436 (
            .O(N__33096),
            .I(N__33093));
    LocalMux I__6435 (
            .O(N__33093),
            .I(N__33090));
    Odrv4 I__6434 (
            .O(N__33090),
            .I(\current_shift_inst.un4_control_input1_1 ));
    InMux I__6433 (
            .O(N__33087),
            .I(N__33083));
    InMux I__6432 (
            .O(N__33086),
            .I(N__33080));
    LocalMux I__6431 (
            .O(N__33083),
            .I(N__33073));
    LocalMux I__6430 (
            .O(N__33080),
            .I(N__33073));
    InMux I__6429 (
            .O(N__33079),
            .I(N__33070));
    InMux I__6428 (
            .O(N__33078),
            .I(N__33067));
    Odrv12 I__6427 (
            .O(N__33073),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6426 (
            .O(N__33070),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6425 (
            .O(N__33067),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__6424 (
            .O(N__33060),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    CascadeMux I__6423 (
            .O(N__33057),
            .I(N__33054));
    InMux I__6422 (
            .O(N__33054),
            .I(N__33051));
    LocalMux I__6421 (
            .O(N__33051),
            .I(N__33048));
    Span4Mux_h I__6420 (
            .O(N__33048),
            .I(N__33045));
    Odrv4 I__6419 (
            .O(N__33045),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    InMux I__6418 (
            .O(N__33042),
            .I(N__33032));
    InMux I__6417 (
            .O(N__33041),
            .I(N__33032));
    InMux I__6416 (
            .O(N__33040),
            .I(N__33032));
    InMux I__6415 (
            .O(N__33039),
            .I(N__33029));
    LocalMux I__6414 (
            .O(N__33032),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__6413 (
            .O(N__33029),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    CascadeMux I__6412 (
            .O(N__33024),
            .I(N__33021));
    InMux I__6411 (
            .O(N__33021),
            .I(N__33013));
    InMux I__6410 (
            .O(N__33020),
            .I(N__33013));
    InMux I__6409 (
            .O(N__33019),
            .I(N__33010));
    InMux I__6408 (
            .O(N__33018),
            .I(N__33007));
    LocalMux I__6407 (
            .O(N__33013),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6406 (
            .O(N__33010),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6405 (
            .O(N__33007),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__6404 (
            .O(N__33000),
            .I(N__32997));
    LocalMux I__6403 (
            .O(N__32997),
            .I(N__32994));
    Odrv12 I__6402 (
            .O(N__32994),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    InMux I__6401 (
            .O(N__32991),
            .I(bfn_13_22_0_));
    InMux I__6400 (
            .O(N__32988),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__6399 (
            .O(N__32985),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__6398 (
            .O(N__32982),
            .I(N__32979));
    LocalMux I__6397 (
            .O(N__32979),
            .I(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ));
    CascadeMux I__6396 (
            .O(N__32976),
            .I(N__32973));
    InMux I__6395 (
            .O(N__32973),
            .I(N__32970));
    LocalMux I__6394 (
            .O(N__32970),
            .I(N__32967));
    Odrv4 I__6393 (
            .O(N__32967),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__6392 (
            .O(N__32964),
            .I(N__32961));
    LocalMux I__6391 (
            .O(N__32961),
            .I(N__32958));
    Span4Mux_h I__6390 (
            .O(N__32958),
            .I(N__32955));
    Odrv4 I__6389 (
            .O(N__32955),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    CascadeMux I__6388 (
            .O(N__32952),
            .I(N__32949));
    InMux I__6387 (
            .O(N__32949),
            .I(N__32946));
    LocalMux I__6386 (
            .O(N__32946),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__6385 (
            .O(N__32943),
            .I(N__32940));
    LocalMux I__6384 (
            .O(N__32940),
            .I(N__32937));
    Odrv4 I__6383 (
            .O(N__32937),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__6382 (
            .O(N__32934),
            .I(N__32931));
    LocalMux I__6381 (
            .O(N__32931),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    CascadeMux I__6380 (
            .O(N__32928),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    InMux I__6379 (
            .O(N__32925),
            .I(N__32922));
    LocalMux I__6378 (
            .O(N__32922),
            .I(N__32918));
    InMux I__6377 (
            .O(N__32921),
            .I(N__32915));
    Odrv12 I__6376 (
            .O(N__32918),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    LocalMux I__6375 (
            .O(N__32915),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    InMux I__6374 (
            .O(N__32910),
            .I(N__32907));
    LocalMux I__6373 (
            .O(N__32907),
            .I(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ));
    InMux I__6372 (
            .O(N__32904),
            .I(N__32901));
    LocalMux I__6371 (
            .O(N__32901),
            .I(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ));
    InMux I__6370 (
            .O(N__32898),
            .I(N__32895));
    LocalMux I__6369 (
            .O(N__32895),
            .I(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ));
    CascadeMux I__6368 (
            .O(N__32892),
            .I(N__32888));
    InMux I__6367 (
            .O(N__32891),
            .I(N__32885));
    InMux I__6366 (
            .O(N__32888),
            .I(N__32882));
    LocalMux I__6365 (
            .O(N__32885),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    LocalMux I__6364 (
            .O(N__32882),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    InMux I__6363 (
            .O(N__32877),
            .I(N__32874));
    LocalMux I__6362 (
            .O(N__32874),
            .I(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ));
    CascadeMux I__6361 (
            .O(N__32871),
            .I(N__32868));
    InMux I__6360 (
            .O(N__32868),
            .I(N__32865));
    LocalMux I__6359 (
            .O(N__32865),
            .I(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ));
    InMux I__6358 (
            .O(N__32862),
            .I(N__32859));
    LocalMux I__6357 (
            .O(N__32859),
            .I(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ));
    CascadeMux I__6356 (
            .O(N__32856),
            .I(N__32853));
    InMux I__6355 (
            .O(N__32853),
            .I(N__32850));
    LocalMux I__6354 (
            .O(N__32850),
            .I(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ));
    InMux I__6353 (
            .O(N__32847),
            .I(N__32844));
    LocalMux I__6352 (
            .O(N__32844),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    CascadeMux I__6351 (
            .O(N__32841),
            .I(N__32838));
    InMux I__6350 (
            .O(N__32838),
            .I(N__32835));
    LocalMux I__6349 (
            .O(N__32835),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    InMux I__6348 (
            .O(N__32832),
            .I(N__32829));
    LocalMux I__6347 (
            .O(N__32829),
            .I(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ));
    CascadeMux I__6346 (
            .O(N__32826),
            .I(N__32823));
    InMux I__6345 (
            .O(N__32823),
            .I(N__32820));
    LocalMux I__6344 (
            .O(N__32820),
            .I(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ));
    CascadeMux I__6343 (
            .O(N__32817),
            .I(N__32814));
    InMux I__6342 (
            .O(N__32814),
            .I(N__32811));
    LocalMux I__6341 (
            .O(N__32811),
            .I(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ));
    CascadeMux I__6340 (
            .O(N__32808),
            .I(N__32804));
    CascadeMux I__6339 (
            .O(N__32807),
            .I(N__32801));
    InMux I__6338 (
            .O(N__32804),
            .I(N__32798));
    InMux I__6337 (
            .O(N__32801),
            .I(N__32793));
    LocalMux I__6336 (
            .O(N__32798),
            .I(N__32790));
    InMux I__6335 (
            .O(N__32797),
            .I(N__32787));
    InMux I__6334 (
            .O(N__32796),
            .I(N__32784));
    LocalMux I__6333 (
            .O(N__32793),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__6332 (
            .O(N__32790),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__6331 (
            .O(N__32787),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__6330 (
            .O(N__32784),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__6329 (
            .O(N__32775),
            .I(N__32772));
    InMux I__6328 (
            .O(N__32772),
            .I(N__32769));
    LocalMux I__6327 (
            .O(N__32769),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__6326 (
            .O(N__32766),
            .I(N__32763));
    LocalMux I__6325 (
            .O(N__32763),
            .I(N__32760));
    Span4Mux_v I__6324 (
            .O(N__32760),
            .I(N__32757));
    Odrv4 I__6323 (
            .O(N__32757),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CascadeMux I__6322 (
            .O(N__32754),
            .I(N__32750));
    CascadeMux I__6321 (
            .O(N__32753),
            .I(N__32746));
    InMux I__6320 (
            .O(N__32750),
            .I(N__32741));
    InMux I__6319 (
            .O(N__32749),
            .I(N__32741));
    InMux I__6318 (
            .O(N__32746),
            .I(N__32738));
    LocalMux I__6317 (
            .O(N__32741),
            .I(N__32735));
    LocalMux I__6316 (
            .O(N__32738),
            .I(N__32732));
    Span4Mux_v I__6315 (
            .O(N__32735),
            .I(N__32726));
    Span4Mux_v I__6314 (
            .O(N__32732),
            .I(N__32726));
    InMux I__6313 (
            .O(N__32731),
            .I(N__32723));
    Span4Mux_v I__6312 (
            .O(N__32726),
            .I(N__32720));
    LocalMux I__6311 (
            .O(N__32723),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__6310 (
            .O(N__32720),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__6309 (
            .O(N__32715),
            .I(N__32710));
    InMux I__6308 (
            .O(N__32714),
            .I(N__32705));
    InMux I__6307 (
            .O(N__32713),
            .I(N__32705));
    LocalMux I__6306 (
            .O(N__32710),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__6305 (
            .O(N__32705),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__6304 (
            .O(N__32700),
            .I(N__32696));
    InMux I__6303 (
            .O(N__32699),
            .I(N__32693));
    LocalMux I__6302 (
            .O(N__32696),
            .I(N__32690));
    LocalMux I__6301 (
            .O(N__32693),
            .I(N__32684));
    Span4Mux_v I__6300 (
            .O(N__32690),
            .I(N__32684));
    InMux I__6299 (
            .O(N__32689),
            .I(N__32681));
    Sp12to4 I__6298 (
            .O(N__32684),
            .I(N__32678));
    LocalMux I__6297 (
            .O(N__32681),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv12 I__6296 (
            .O(N__32678),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__6295 (
            .O(N__32673),
            .I(N__32669));
    InMux I__6294 (
            .O(N__32672),
            .I(N__32666));
    LocalMux I__6293 (
            .O(N__32669),
            .I(N__32661));
    LocalMux I__6292 (
            .O(N__32666),
            .I(N__32661));
    Span4Mux_s3_v I__6291 (
            .O(N__32661),
            .I(N__32658));
    Span4Mux_h I__6290 (
            .O(N__32658),
            .I(N__32655));
    Sp12to4 I__6289 (
            .O(N__32655),
            .I(N__32650));
    InMux I__6288 (
            .O(N__32654),
            .I(N__32645));
    InMux I__6287 (
            .O(N__32653),
            .I(N__32645));
    Span12Mux_v I__6286 (
            .O(N__32650),
            .I(N__32642));
    LocalMux I__6285 (
            .O(N__32645),
            .I(N__32639));
    Span12Mux_v I__6284 (
            .O(N__32642),
            .I(N__32636));
    Span12Mux_h I__6283 (
            .O(N__32639),
            .I(N__32633));
    Span12Mux_h I__6282 (
            .O(N__32636),
            .I(N__32628));
    Span12Mux_v I__6281 (
            .O(N__32633),
            .I(N__32628));
    Odrv12 I__6280 (
            .O(N__32628),
            .I(start_stop_c));
    InMux I__6279 (
            .O(N__32625),
            .I(N__32622));
    LocalMux I__6278 (
            .O(N__32622),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    CascadeMux I__6277 (
            .O(N__32619),
            .I(N__32616));
    InMux I__6276 (
            .O(N__32616),
            .I(N__32610));
    InMux I__6275 (
            .O(N__32615),
            .I(N__32610));
    LocalMux I__6274 (
            .O(N__32610),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    CascadeMux I__6273 (
            .O(N__32607),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_));
    InMux I__6272 (
            .O(N__32604),
            .I(N__32598));
    InMux I__6271 (
            .O(N__32603),
            .I(N__32598));
    LocalMux I__6270 (
            .O(N__32598),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ));
    CascadeMux I__6269 (
            .O(N__32595),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_));
    InMux I__6268 (
            .O(N__32592),
            .I(N__32583));
    InMux I__6267 (
            .O(N__32591),
            .I(N__32583));
    InMux I__6266 (
            .O(N__32590),
            .I(N__32583));
    LocalMux I__6265 (
            .O(N__32583),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    InMux I__6264 (
            .O(N__32580),
            .I(N__32571));
    InMux I__6263 (
            .O(N__32579),
            .I(N__32571));
    InMux I__6262 (
            .O(N__32578),
            .I(N__32571));
    LocalMux I__6261 (
            .O(N__32571),
            .I(N__32568));
    Span4Mux_v I__6260 (
            .O(N__32568),
            .I(N__32565));
    Odrv4 I__6259 (
            .O(N__32565),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    InMux I__6258 (
            .O(N__32562),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__6257 (
            .O(N__32559),
            .I(bfn_13_10_0_));
    InMux I__6256 (
            .O(N__32556),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__6255 (
            .O(N__32553),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__6254 (
            .O(N__32550),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__6253 (
            .O(N__32547),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__6252 (
            .O(N__32544),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23_cascade_));
    InMux I__6251 (
            .O(N__32541),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__6250 (
            .O(N__32538),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__6249 (
            .O(N__32535),
            .I(bfn_13_9_0_));
    InMux I__6248 (
            .O(N__32532),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__6247 (
            .O(N__32529),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__6246 (
            .O(N__32526),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__6245 (
            .O(N__32523),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__6244 (
            .O(N__32520),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__6243 (
            .O(N__32517),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__6242 (
            .O(N__32514),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__6241 (
            .O(N__32511),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__6240 (
            .O(N__32508),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__6239 (
            .O(N__32505),
            .I(bfn_13_8_0_));
    InMux I__6238 (
            .O(N__32502),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__6237 (
            .O(N__32499),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__6236 (
            .O(N__32496),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__6235 (
            .O(N__32493),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__6234 (
            .O(N__32490),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    IoInMux I__6233 (
            .O(N__32487),
            .I(N__32484));
    LocalMux I__6232 (
            .O(N__32484),
            .I(N__32481));
    Span4Mux_s0_v I__6231 (
            .O(N__32481),
            .I(N__32471));
    InMux I__6230 (
            .O(N__32480),
            .I(N__32440));
    InMux I__6229 (
            .O(N__32479),
            .I(N__32440));
    InMux I__6228 (
            .O(N__32478),
            .I(N__32440));
    InMux I__6227 (
            .O(N__32477),
            .I(N__32431));
    InMux I__6226 (
            .O(N__32476),
            .I(N__32431));
    InMux I__6225 (
            .O(N__32475),
            .I(N__32431));
    InMux I__6224 (
            .O(N__32474),
            .I(N__32431));
    Sp12to4 I__6223 (
            .O(N__32471),
            .I(N__32428));
    InMux I__6222 (
            .O(N__32470),
            .I(N__32425));
    InMux I__6221 (
            .O(N__32469),
            .I(N__32416));
    InMux I__6220 (
            .O(N__32468),
            .I(N__32416));
    InMux I__6219 (
            .O(N__32467),
            .I(N__32416));
    InMux I__6218 (
            .O(N__32466),
            .I(N__32416));
    InMux I__6217 (
            .O(N__32465),
            .I(N__32407));
    InMux I__6216 (
            .O(N__32464),
            .I(N__32407));
    InMux I__6215 (
            .O(N__32463),
            .I(N__32407));
    InMux I__6214 (
            .O(N__32462),
            .I(N__32407));
    InMux I__6213 (
            .O(N__32461),
            .I(N__32400));
    InMux I__6212 (
            .O(N__32460),
            .I(N__32400));
    InMux I__6211 (
            .O(N__32459),
            .I(N__32400));
    InMux I__6210 (
            .O(N__32458),
            .I(N__32391));
    InMux I__6209 (
            .O(N__32457),
            .I(N__32391));
    InMux I__6208 (
            .O(N__32456),
            .I(N__32391));
    InMux I__6207 (
            .O(N__32455),
            .I(N__32391));
    InMux I__6206 (
            .O(N__32454),
            .I(N__32382));
    InMux I__6205 (
            .O(N__32453),
            .I(N__32382));
    InMux I__6204 (
            .O(N__32452),
            .I(N__32382));
    InMux I__6203 (
            .O(N__32451),
            .I(N__32382));
    InMux I__6202 (
            .O(N__32450),
            .I(N__32373));
    InMux I__6201 (
            .O(N__32449),
            .I(N__32373));
    InMux I__6200 (
            .O(N__32448),
            .I(N__32373));
    InMux I__6199 (
            .O(N__32447),
            .I(N__32373));
    LocalMux I__6198 (
            .O(N__32440),
            .I(N__32368));
    LocalMux I__6197 (
            .O(N__32431),
            .I(N__32368));
    Span12Mux_s5_h I__6196 (
            .O(N__32428),
            .I(N__32365));
    LocalMux I__6195 (
            .O(N__32425),
            .I(N__32362));
    LocalMux I__6194 (
            .O(N__32416),
            .I(N__32357));
    LocalMux I__6193 (
            .O(N__32407),
            .I(N__32357));
    LocalMux I__6192 (
            .O(N__32400),
            .I(N__32348));
    LocalMux I__6191 (
            .O(N__32391),
            .I(N__32348));
    LocalMux I__6190 (
            .O(N__32382),
            .I(N__32348));
    LocalMux I__6189 (
            .O(N__32373),
            .I(N__32348));
    Span4Mux_h I__6188 (
            .O(N__32368),
            .I(N__32345));
    Span12Mux_v I__6187 (
            .O(N__32365),
            .I(N__32342));
    Span12Mux_h I__6186 (
            .O(N__32362),
            .I(N__32339));
    Span4Mux_v I__6185 (
            .O(N__32357),
            .I(N__32334));
    Span4Mux_v I__6184 (
            .O(N__32348),
            .I(N__32334));
    Span4Mux_v I__6183 (
            .O(N__32345),
            .I(N__32331));
    Span12Mux_v I__6182 (
            .O(N__32342),
            .I(N__32328));
    Odrv12 I__6181 (
            .O(N__32339),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__6180 (
            .O(N__32334),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__6179 (
            .O(N__32331),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__6178 (
            .O(N__32328),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__6177 (
            .O(N__32319),
            .I(N__32316));
    LocalMux I__6176 (
            .O(N__32316),
            .I(N__32312));
    CascadeMux I__6175 (
            .O(N__32315),
            .I(N__32309));
    Span4Mux_h I__6174 (
            .O(N__32312),
            .I(N__32306));
    InMux I__6173 (
            .O(N__32309),
            .I(N__32303));
    Span4Mux_v I__6172 (
            .O(N__32306),
            .I(N__32300));
    LocalMux I__6171 (
            .O(N__32303),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    Odrv4 I__6170 (
            .O(N__32300),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    CascadeMux I__6169 (
            .O(N__32295),
            .I(N__32291));
    InMux I__6168 (
            .O(N__32294),
            .I(N__32280));
    InMux I__6167 (
            .O(N__32291),
            .I(N__32280));
    InMux I__6166 (
            .O(N__32290),
            .I(N__32280));
    InMux I__6165 (
            .O(N__32289),
            .I(N__32280));
    LocalMux I__6164 (
            .O(N__32280),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__6163 (
            .O(N__32277),
            .I(N__32265));
    InMux I__6162 (
            .O(N__32276),
            .I(N__32265));
    InMux I__6161 (
            .O(N__32275),
            .I(N__32265));
    InMux I__6160 (
            .O(N__32274),
            .I(N__32265));
    LocalMux I__6159 (
            .O(N__32265),
            .I(N__32262));
    Span4Mux_v I__6158 (
            .O(N__32262),
            .I(N__32259));
    Odrv4 I__6157 (
            .O(N__32259),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__6156 (
            .O(N__32256),
            .I(N__32253));
    LocalMux I__6155 (
            .O(N__32253),
            .I(N__32250));
    Span4Mux_h I__6154 (
            .O(N__32250),
            .I(N__32246));
    InMux I__6153 (
            .O(N__32249),
            .I(N__32243));
    Span4Mux_v I__6152 (
            .O(N__32246),
            .I(N__32240));
    LocalMux I__6151 (
            .O(N__32243),
            .I(N__32237));
    Odrv4 I__6150 (
            .O(N__32240),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv12 I__6149 (
            .O(N__32237),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    CascadeMux I__6148 (
            .O(N__32232),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ));
    InMux I__6147 (
            .O(N__32229),
            .I(N__32225));
    InMux I__6146 (
            .O(N__32228),
            .I(N__32222));
    LocalMux I__6145 (
            .O(N__32225),
            .I(N__32217));
    LocalMux I__6144 (
            .O(N__32222),
            .I(N__32217));
    Span4Mux_v I__6143 (
            .O(N__32217),
            .I(N__32211));
    InMux I__6142 (
            .O(N__32216),
            .I(N__32204));
    InMux I__6141 (
            .O(N__32215),
            .I(N__32204));
    InMux I__6140 (
            .O(N__32214),
            .I(N__32204));
    Odrv4 I__6139 (
            .O(N__32211),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__6138 (
            .O(N__32204),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    InMux I__6137 (
            .O(N__32199),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__6136 (
            .O(N__32196),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__6135 (
            .O(N__32193),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__6134 (
            .O(N__32190),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__6133 (
            .O(N__32187),
            .I(N__32184));
    LocalMux I__6132 (
            .O(N__32184),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ));
    CascadeMux I__6131 (
            .O(N__32181),
            .I(N__32178));
    InMux I__6130 (
            .O(N__32178),
            .I(N__32175));
    LocalMux I__6129 (
            .O(N__32175),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ));
    IoInMux I__6128 (
            .O(N__32172),
            .I(N__32169));
    LocalMux I__6127 (
            .O(N__32169),
            .I(N__32166));
    Span4Mux_s0_v I__6126 (
            .O(N__32166),
            .I(N__32163));
    Odrv4 I__6125 (
            .O(N__32163),
            .I(\pll_inst.red_c_i ));
    InMux I__6124 (
            .O(N__32160),
            .I(N__32154));
    InMux I__6123 (
            .O(N__32159),
            .I(N__32147));
    InMux I__6122 (
            .O(N__32158),
            .I(N__32147));
    InMux I__6121 (
            .O(N__32157),
            .I(N__32147));
    LocalMux I__6120 (
            .O(N__32154),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__6119 (
            .O(N__32147),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__6118 (
            .O(N__32142),
            .I(N__32139));
    InMux I__6117 (
            .O(N__32139),
            .I(N__32134));
    InMux I__6116 (
            .O(N__32138),
            .I(N__32129));
    InMux I__6115 (
            .O(N__32137),
            .I(N__32129));
    LocalMux I__6114 (
            .O(N__32134),
            .I(N__32126));
    LocalMux I__6113 (
            .O(N__32129),
            .I(N__32123));
    Span4Mux_h I__6112 (
            .O(N__32126),
            .I(N__32120));
    Span4Mux_v I__6111 (
            .O(N__32123),
            .I(N__32117));
    Odrv4 I__6110 (
            .O(N__32120),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    Odrv4 I__6109 (
            .O(N__32117),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    CEMux I__6108 (
            .O(N__32112),
            .I(N__32108));
    CEMux I__6107 (
            .O(N__32111),
            .I(N__32102));
    LocalMux I__6106 (
            .O(N__32108),
            .I(N__32097));
    CEMux I__6105 (
            .O(N__32107),
            .I(N__32094));
    CEMux I__6104 (
            .O(N__32106),
            .I(N__32091));
    CEMux I__6103 (
            .O(N__32105),
            .I(N__32088));
    LocalMux I__6102 (
            .O(N__32102),
            .I(N__32085));
    CEMux I__6101 (
            .O(N__32101),
            .I(N__32075));
    CEMux I__6100 (
            .O(N__32100),
            .I(N__32072));
    Span4Mux_h I__6099 (
            .O(N__32097),
            .I(N__32062));
    LocalMux I__6098 (
            .O(N__32094),
            .I(N__32062));
    LocalMux I__6097 (
            .O(N__32091),
            .I(N__32057));
    LocalMux I__6096 (
            .O(N__32088),
            .I(N__32057));
    Span4Mux_h I__6095 (
            .O(N__32085),
            .I(N__32054));
    InMux I__6094 (
            .O(N__32084),
            .I(N__32042));
    InMux I__6093 (
            .O(N__32083),
            .I(N__32042));
    InMux I__6092 (
            .O(N__32082),
            .I(N__32042));
    CEMux I__6091 (
            .O(N__32081),
            .I(N__32039));
    CEMux I__6090 (
            .O(N__32080),
            .I(N__32036));
    CEMux I__6089 (
            .O(N__32079),
            .I(N__32033));
    CEMux I__6088 (
            .O(N__32078),
            .I(N__32030));
    LocalMux I__6087 (
            .O(N__32075),
            .I(N__32022));
    LocalMux I__6086 (
            .O(N__32072),
            .I(N__32019));
    CEMux I__6085 (
            .O(N__32071),
            .I(N__32011));
    CEMux I__6084 (
            .O(N__32070),
            .I(N__32008));
    InMux I__6083 (
            .O(N__32069),
            .I(N__32001));
    InMux I__6082 (
            .O(N__32068),
            .I(N__32001));
    InMux I__6081 (
            .O(N__32067),
            .I(N__32001));
    Span4Mux_h I__6080 (
            .O(N__32062),
            .I(N__31994));
    Span4Mux_v I__6079 (
            .O(N__32057),
            .I(N__31994));
    Span4Mux_v I__6078 (
            .O(N__32054),
            .I(N__31994));
    InMux I__6077 (
            .O(N__32053),
            .I(N__31985));
    InMux I__6076 (
            .O(N__32052),
            .I(N__31985));
    InMux I__6075 (
            .O(N__32051),
            .I(N__31985));
    InMux I__6074 (
            .O(N__32050),
            .I(N__31985));
    CEMux I__6073 (
            .O(N__32049),
            .I(N__31981));
    LocalMux I__6072 (
            .O(N__32042),
            .I(N__31978));
    LocalMux I__6071 (
            .O(N__32039),
            .I(N__31975));
    LocalMux I__6070 (
            .O(N__32036),
            .I(N__31968));
    LocalMux I__6069 (
            .O(N__32033),
            .I(N__31968));
    LocalMux I__6068 (
            .O(N__32030),
            .I(N__31968));
    CEMux I__6067 (
            .O(N__32029),
            .I(N__31953));
    InMux I__6066 (
            .O(N__32028),
            .I(N__31944));
    InMux I__6065 (
            .O(N__32027),
            .I(N__31944));
    InMux I__6064 (
            .O(N__32026),
            .I(N__31944));
    InMux I__6063 (
            .O(N__32025),
            .I(N__31944));
    Span4Mux_v I__6062 (
            .O(N__32022),
            .I(N__31939));
    Span4Mux_h I__6061 (
            .O(N__32019),
            .I(N__31939));
    CEMux I__6060 (
            .O(N__32018),
            .I(N__31936));
    InMux I__6059 (
            .O(N__32017),
            .I(N__31927));
    InMux I__6058 (
            .O(N__32016),
            .I(N__31927));
    InMux I__6057 (
            .O(N__32015),
            .I(N__31927));
    InMux I__6056 (
            .O(N__32014),
            .I(N__31927));
    LocalMux I__6055 (
            .O(N__32011),
            .I(N__31924));
    LocalMux I__6054 (
            .O(N__32008),
            .I(N__31921));
    LocalMux I__6053 (
            .O(N__32001),
            .I(N__31918));
    Span4Mux_v I__6052 (
            .O(N__31994),
            .I(N__31913));
    LocalMux I__6051 (
            .O(N__31985),
            .I(N__31913));
    InMux I__6050 (
            .O(N__31984),
            .I(N__31910));
    LocalMux I__6049 (
            .O(N__31981),
            .I(N__31907));
    Span4Mux_h I__6048 (
            .O(N__31978),
            .I(N__31902));
    Span4Mux_h I__6047 (
            .O(N__31975),
            .I(N__31902));
    Span4Mux_v I__6046 (
            .O(N__31968),
            .I(N__31899));
    InMux I__6045 (
            .O(N__31967),
            .I(N__31890));
    InMux I__6044 (
            .O(N__31966),
            .I(N__31890));
    InMux I__6043 (
            .O(N__31965),
            .I(N__31890));
    InMux I__6042 (
            .O(N__31964),
            .I(N__31890));
    InMux I__6041 (
            .O(N__31963),
            .I(N__31881));
    InMux I__6040 (
            .O(N__31962),
            .I(N__31881));
    InMux I__6039 (
            .O(N__31961),
            .I(N__31881));
    InMux I__6038 (
            .O(N__31960),
            .I(N__31881));
    InMux I__6037 (
            .O(N__31959),
            .I(N__31872));
    InMux I__6036 (
            .O(N__31958),
            .I(N__31872));
    InMux I__6035 (
            .O(N__31957),
            .I(N__31872));
    InMux I__6034 (
            .O(N__31956),
            .I(N__31872));
    LocalMux I__6033 (
            .O(N__31953),
            .I(N__31865));
    LocalMux I__6032 (
            .O(N__31944),
            .I(N__31865));
    Span4Mux_h I__6031 (
            .O(N__31939),
            .I(N__31865));
    LocalMux I__6030 (
            .O(N__31936),
            .I(N__31856));
    LocalMux I__6029 (
            .O(N__31927),
            .I(N__31856));
    Span4Mux_v I__6028 (
            .O(N__31924),
            .I(N__31856));
    Span4Mux_v I__6027 (
            .O(N__31921),
            .I(N__31856));
    Span4Mux_h I__6026 (
            .O(N__31918),
            .I(N__31851));
    Span4Mux_h I__6025 (
            .O(N__31913),
            .I(N__31851));
    LocalMux I__6024 (
            .O(N__31910),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv12 I__6023 (
            .O(N__31907),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__6022 (
            .O(N__31902),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__6021 (
            .O(N__31899),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__6020 (
            .O(N__31890),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__6019 (
            .O(N__31881),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__6018 (
            .O(N__31872),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__6017 (
            .O(N__31865),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__6016 (
            .O(N__31856),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__6015 (
            .O(N__31851),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__6014 (
            .O(N__31830),
            .I(N__31827));
    LocalMux I__6013 (
            .O(N__31827),
            .I(N__31823));
    InMux I__6012 (
            .O(N__31826),
            .I(N__31819));
    Span4Mux_h I__6011 (
            .O(N__31823),
            .I(N__31816));
    InMux I__6010 (
            .O(N__31822),
            .I(N__31813));
    LocalMux I__6009 (
            .O(N__31819),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__6008 (
            .O(N__31816),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__6007 (
            .O(N__31813),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__6006 (
            .O(N__31806),
            .I(N__31803));
    LocalMux I__6005 (
            .O(N__31803),
            .I(N__31800));
    Odrv4 I__6004 (
            .O(N__31800),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    IoInMux I__6003 (
            .O(N__31797),
            .I(N__31794));
    LocalMux I__6002 (
            .O(N__31794),
            .I(N__31791));
    Span4Mux_s2_v I__6001 (
            .O(N__31791),
            .I(N__31788));
    Span4Mux_h I__6000 (
            .O(N__31788),
            .I(N__31785));
    Span4Mux_v I__5999 (
            .O(N__31785),
            .I(N__31780));
    InMux I__5998 (
            .O(N__31784),
            .I(N__31775));
    InMux I__5997 (
            .O(N__31783),
            .I(N__31775));
    Odrv4 I__5996 (
            .O(N__31780),
            .I(s1_phy_c));
    LocalMux I__5995 (
            .O(N__31775),
            .I(s1_phy_c));
    InMux I__5994 (
            .O(N__31770),
            .I(N__31761));
    InMux I__5993 (
            .O(N__31769),
            .I(N__31761));
    InMux I__5992 (
            .O(N__31768),
            .I(N__31761));
    LocalMux I__5991 (
            .O(N__31761),
            .I(N__31756));
    InMux I__5990 (
            .O(N__31760),
            .I(N__31752));
    InMux I__5989 (
            .O(N__31759),
            .I(N__31749));
    Span4Mux_v I__5988 (
            .O(N__31756),
            .I(N__31746));
    InMux I__5987 (
            .O(N__31755),
            .I(N__31743));
    LocalMux I__5986 (
            .O(N__31752),
            .I(state_3));
    LocalMux I__5985 (
            .O(N__31749),
            .I(state_3));
    Odrv4 I__5984 (
            .O(N__31746),
            .I(state_3));
    LocalMux I__5983 (
            .O(N__31743),
            .I(state_3));
    InMux I__5982 (
            .O(N__31734),
            .I(N__31731));
    LocalMux I__5981 (
            .O(N__31731),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ));
    CascadeMux I__5980 (
            .O(N__31728),
            .I(N__31725));
    InMux I__5979 (
            .O(N__31725),
            .I(N__31722));
    LocalMux I__5978 (
            .O(N__31722),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ));
    InMux I__5977 (
            .O(N__31719),
            .I(N__31716));
    LocalMux I__5976 (
            .O(N__31716),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ));
    CascadeMux I__5975 (
            .O(N__31713),
            .I(N__31710));
    InMux I__5974 (
            .O(N__31710),
            .I(N__31707));
    LocalMux I__5973 (
            .O(N__31707),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ));
    CascadeMux I__5972 (
            .O(N__31704),
            .I(N__31701));
    InMux I__5971 (
            .O(N__31701),
            .I(N__31698));
    LocalMux I__5970 (
            .O(N__31698),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ));
    InMux I__5969 (
            .O(N__31695),
            .I(N__31692));
    LocalMux I__5968 (
            .O(N__31692),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ));
    CascadeMux I__5967 (
            .O(N__31689),
            .I(N__31686));
    InMux I__5966 (
            .O(N__31686),
            .I(N__31683));
    LocalMux I__5965 (
            .O(N__31683),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ));
    InMux I__5964 (
            .O(N__31680),
            .I(N__31677));
    LocalMux I__5963 (
            .O(N__31677),
            .I(N__31674));
    Span4Mux_h I__5962 (
            .O(N__31674),
            .I(N__31671));
    Odrv4 I__5961 (
            .O(N__31671),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__5960 (
            .O(N__31668),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    CascadeMux I__5959 (
            .O(N__31665),
            .I(N__31662));
    InMux I__5958 (
            .O(N__31662),
            .I(N__31659));
    LocalMux I__5957 (
            .O(N__31659),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__5956 (
            .O(N__31656),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__5955 (
            .O(N__31653),
            .I(N__31650));
    LocalMux I__5954 (
            .O(N__31650),
            .I(N__31647));
    Span4Mux_h I__5953 (
            .O(N__31647),
            .I(N__31644));
    Odrv4 I__5952 (
            .O(N__31644),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__5951 (
            .O(N__31641),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__5950 (
            .O(N__31638),
            .I(N__31635));
    LocalMux I__5949 (
            .O(N__31635),
            .I(N__31632));
    Odrv4 I__5948 (
            .O(N__31632),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__5947 (
            .O(N__31629),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__5946 (
            .O(N__31626),
            .I(N__31623));
    LocalMux I__5945 (
            .O(N__31623),
            .I(N__31620));
    Odrv4 I__5944 (
            .O(N__31620),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__5943 (
            .O(N__31617),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__5942 (
            .O(N__31614),
            .I(N__31611));
    LocalMux I__5941 (
            .O(N__31611),
            .I(N__31608));
    Odrv4 I__5940 (
            .O(N__31608),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__5939 (
            .O(N__31605),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__5938 (
            .O(N__31602),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__5937 (
            .O(N__31599),
            .I(N__31596));
    LocalMux I__5936 (
            .O(N__31596),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__5935 (
            .O(N__31593),
            .I(N__31590));
    LocalMux I__5934 (
            .O(N__31590),
            .I(N__31587));
    Span4Mux_v I__5933 (
            .O(N__31587),
            .I(N__31584));
    Odrv4 I__5932 (
            .O(N__31584),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__5931 (
            .O(N__31581),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__5930 (
            .O(N__31578),
            .I(N__31575));
    LocalMux I__5929 (
            .O(N__31575),
            .I(N__31572));
    Span4Mux_v I__5928 (
            .O(N__31572),
            .I(N__31569));
    Odrv4 I__5927 (
            .O(N__31569),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__5926 (
            .O(N__31566),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__5925 (
            .O(N__31563),
            .I(N__31560));
    LocalMux I__5924 (
            .O(N__31560),
            .I(N__31557));
    Span4Mux_h I__5923 (
            .O(N__31557),
            .I(N__31554));
    Odrv4 I__5922 (
            .O(N__31554),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__5921 (
            .O(N__31551),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__5920 (
            .O(N__31548),
            .I(N__31545));
    LocalMux I__5919 (
            .O(N__31545),
            .I(N__31542));
    Span4Mux_h I__5918 (
            .O(N__31542),
            .I(N__31539));
    Odrv4 I__5917 (
            .O(N__31539),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__5916 (
            .O(N__31536),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__5915 (
            .O(N__31533),
            .I(N__31530));
    LocalMux I__5914 (
            .O(N__31530),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__5913 (
            .O(N__31527),
            .I(bfn_12_20_0_));
    CascadeMux I__5912 (
            .O(N__31524),
            .I(N__31521));
    InMux I__5911 (
            .O(N__31521),
            .I(N__31518));
    LocalMux I__5910 (
            .O(N__31518),
            .I(N__31515));
    Odrv12 I__5909 (
            .O(N__31515),
            .I(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ));
    CascadeMux I__5908 (
            .O(N__31512),
            .I(N__31509));
    InMux I__5907 (
            .O(N__31509),
            .I(N__31506));
    LocalMux I__5906 (
            .O(N__31506),
            .I(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ));
    CascadeMux I__5905 (
            .O(N__31503),
            .I(N__31500));
    InMux I__5904 (
            .O(N__31500),
            .I(N__31497));
    LocalMux I__5903 (
            .O(N__31497),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    InMux I__5902 (
            .O(N__31494),
            .I(N__31484));
    InMux I__5901 (
            .O(N__31493),
            .I(N__31484));
    InMux I__5900 (
            .O(N__31492),
            .I(N__31484));
    InMux I__5899 (
            .O(N__31491),
            .I(N__31481));
    LocalMux I__5898 (
            .O(N__31484),
            .I(N__31478));
    LocalMux I__5897 (
            .O(N__31481),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__5896 (
            .O(N__31478),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__5895 (
            .O(N__31473),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__5894 (
            .O(N__31470),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    CascadeMux I__5893 (
            .O(N__31467),
            .I(N__31463));
    CascadeMux I__5892 (
            .O(N__31466),
            .I(N__31459));
    InMux I__5891 (
            .O(N__31463),
            .I(N__31452));
    InMux I__5890 (
            .O(N__31462),
            .I(N__31452));
    InMux I__5889 (
            .O(N__31459),
            .I(N__31452));
    LocalMux I__5888 (
            .O(N__31452),
            .I(N__31448));
    InMux I__5887 (
            .O(N__31451),
            .I(N__31445));
    Span4Mux_h I__5886 (
            .O(N__31448),
            .I(N__31442));
    LocalMux I__5885 (
            .O(N__31445),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__5884 (
            .O(N__31442),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__5883 (
            .O(N__31437),
            .I(N__31433));
    InMux I__5882 (
            .O(N__31436),
            .I(N__31429));
    InMux I__5881 (
            .O(N__31433),
            .I(N__31426));
    InMux I__5880 (
            .O(N__31432),
            .I(N__31423));
    LocalMux I__5879 (
            .O(N__31429),
            .I(il_max_comp1_D2));
    LocalMux I__5878 (
            .O(N__31426),
            .I(il_max_comp1_D2));
    LocalMux I__5877 (
            .O(N__31423),
            .I(il_max_comp1_D2));
    CascadeMux I__5876 (
            .O(N__31416),
            .I(N__31413));
    InMux I__5875 (
            .O(N__31413),
            .I(N__31410));
    LocalMux I__5874 (
            .O(N__31410),
            .I(N__31407));
    Odrv4 I__5873 (
            .O(N__31407),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    InMux I__5872 (
            .O(N__31404),
            .I(N__31401));
    LocalMux I__5871 (
            .O(N__31401),
            .I(N__31398));
    Odrv4 I__5870 (
            .O(N__31398),
            .I(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ));
    CascadeMux I__5869 (
            .O(N__31395),
            .I(N__31392));
    InMux I__5868 (
            .O(N__31392),
            .I(N__31389));
    LocalMux I__5867 (
            .O(N__31389),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    CascadeMux I__5866 (
            .O(N__31386),
            .I(N__31383));
    InMux I__5865 (
            .O(N__31383),
            .I(N__31380));
    LocalMux I__5864 (
            .O(N__31380),
            .I(N__31377));
    Odrv4 I__5863 (
            .O(N__31377),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ));
    CascadeMux I__5862 (
            .O(N__31374),
            .I(N__31371));
    InMux I__5861 (
            .O(N__31371),
            .I(N__31365));
    InMux I__5860 (
            .O(N__31370),
            .I(N__31365));
    LocalMux I__5859 (
            .O(N__31365),
            .I(N__31361));
    InMux I__5858 (
            .O(N__31364),
            .I(N__31358));
    Span4Mux_h I__5857 (
            .O(N__31361),
            .I(N__31355));
    LocalMux I__5856 (
            .O(N__31358),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__5855 (
            .O(N__31355),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__5854 (
            .O(N__31350),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__5853 (
            .O(N__31347),
            .I(N__31341));
    InMux I__5852 (
            .O(N__31346),
            .I(N__31341));
    LocalMux I__5851 (
            .O(N__31341),
            .I(N__31337));
    InMux I__5850 (
            .O(N__31340),
            .I(N__31334));
    Span4Mux_h I__5849 (
            .O(N__31337),
            .I(N__31331));
    LocalMux I__5848 (
            .O(N__31334),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__5847 (
            .O(N__31331),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__5846 (
            .O(N__31326),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    CascadeMux I__5845 (
            .O(N__31323),
            .I(N__31320));
    InMux I__5844 (
            .O(N__31320),
            .I(N__31314));
    InMux I__5843 (
            .O(N__31319),
            .I(N__31314));
    LocalMux I__5842 (
            .O(N__31314),
            .I(N__31310));
    InMux I__5841 (
            .O(N__31313),
            .I(N__31307));
    Span4Mux_h I__5840 (
            .O(N__31310),
            .I(N__31304));
    LocalMux I__5839 (
            .O(N__31307),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__5838 (
            .O(N__31304),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__5837 (
            .O(N__31299),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__5836 (
            .O(N__31296),
            .I(N__31289));
    InMux I__5835 (
            .O(N__31295),
            .I(N__31289));
    InMux I__5834 (
            .O(N__31294),
            .I(N__31286));
    LocalMux I__5833 (
            .O(N__31289),
            .I(N__31283));
    LocalMux I__5832 (
            .O(N__31286),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__5831 (
            .O(N__31283),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__5830 (
            .O(N__31278),
            .I(bfn_12_13_0_));
    InMux I__5829 (
            .O(N__31275),
            .I(N__31271));
    CascadeMux I__5828 (
            .O(N__31274),
            .I(N__31268));
    LocalMux I__5827 (
            .O(N__31271),
            .I(N__31264));
    InMux I__5826 (
            .O(N__31268),
            .I(N__31261));
    InMux I__5825 (
            .O(N__31267),
            .I(N__31258));
    Span4Mux_v I__5824 (
            .O(N__31264),
            .I(N__31253));
    LocalMux I__5823 (
            .O(N__31261),
            .I(N__31253));
    LocalMux I__5822 (
            .O(N__31258),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    Odrv4 I__5821 (
            .O(N__31253),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__5820 (
            .O(N__31248),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    CascadeMux I__5819 (
            .O(N__31245),
            .I(N__31242));
    InMux I__5818 (
            .O(N__31242),
            .I(N__31238));
    InMux I__5817 (
            .O(N__31241),
            .I(N__31234));
    LocalMux I__5816 (
            .O(N__31238),
            .I(N__31231));
    InMux I__5815 (
            .O(N__31237),
            .I(N__31228));
    LocalMux I__5814 (
            .O(N__31234),
            .I(N__31225));
    Span4Mux_h I__5813 (
            .O(N__31231),
            .I(N__31222));
    LocalMux I__5812 (
            .O(N__31228),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv4 I__5811 (
            .O(N__31225),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv4 I__5810 (
            .O(N__31222),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__5809 (
            .O(N__31215),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    CascadeMux I__5808 (
            .O(N__31212),
            .I(N__31209));
    InMux I__5807 (
            .O(N__31209),
            .I(N__31203));
    InMux I__5806 (
            .O(N__31208),
            .I(N__31203));
    LocalMux I__5805 (
            .O(N__31203),
            .I(N__31199));
    InMux I__5804 (
            .O(N__31202),
            .I(N__31196));
    Span4Mux_h I__5803 (
            .O(N__31199),
            .I(N__31193));
    LocalMux I__5802 (
            .O(N__31196),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv4 I__5801 (
            .O(N__31193),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__5800 (
            .O(N__31188),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__5799 (
            .O(N__31185),
            .I(N__31179));
    InMux I__5798 (
            .O(N__31184),
            .I(N__31179));
    LocalMux I__5797 (
            .O(N__31179),
            .I(N__31175));
    InMux I__5796 (
            .O(N__31178),
            .I(N__31172));
    Span4Mux_h I__5795 (
            .O(N__31175),
            .I(N__31169));
    LocalMux I__5794 (
            .O(N__31172),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__5793 (
            .O(N__31169),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__5792 (
            .O(N__31164),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__5791 (
            .O(N__31161),
            .I(N__31157));
    InMux I__5790 (
            .O(N__31160),
            .I(N__31154));
    LocalMux I__5789 (
            .O(N__31157),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__5788 (
            .O(N__31154),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__5787 (
            .O(N__31149),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__5786 (
            .O(N__31146),
            .I(N__31142));
    InMux I__5785 (
            .O(N__31145),
            .I(N__31139));
    LocalMux I__5784 (
            .O(N__31142),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__5783 (
            .O(N__31139),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__5782 (
            .O(N__31134),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__5781 (
            .O(N__31131),
            .I(N__31127));
    InMux I__5780 (
            .O(N__31130),
            .I(N__31124));
    LocalMux I__5779 (
            .O(N__31127),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__5778 (
            .O(N__31124),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__5777 (
            .O(N__31119),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    CascadeMux I__5776 (
            .O(N__31116),
            .I(N__31113));
    InMux I__5775 (
            .O(N__31113),
            .I(N__31107));
    InMux I__5774 (
            .O(N__31112),
            .I(N__31107));
    LocalMux I__5773 (
            .O(N__31107),
            .I(N__31103));
    InMux I__5772 (
            .O(N__31106),
            .I(N__31100));
    Span4Mux_h I__5771 (
            .O(N__31103),
            .I(N__31097));
    LocalMux I__5770 (
            .O(N__31100),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__5769 (
            .O(N__31097),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__5768 (
            .O(N__31092),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__5767 (
            .O(N__31089),
            .I(N__31082));
    InMux I__5766 (
            .O(N__31088),
            .I(N__31082));
    InMux I__5765 (
            .O(N__31087),
            .I(N__31079));
    LocalMux I__5764 (
            .O(N__31082),
            .I(N__31076));
    LocalMux I__5763 (
            .O(N__31079),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv12 I__5762 (
            .O(N__31076),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__5761 (
            .O(N__31071),
            .I(bfn_12_12_0_));
    InMux I__5760 (
            .O(N__31068),
            .I(N__31062));
    InMux I__5759 (
            .O(N__31067),
            .I(N__31062));
    LocalMux I__5758 (
            .O(N__31062),
            .I(N__31058));
    InMux I__5757 (
            .O(N__31061),
            .I(N__31055));
    Span4Mux_h I__5756 (
            .O(N__31058),
            .I(N__31052));
    LocalMux I__5755 (
            .O(N__31055),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__5754 (
            .O(N__31052),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__5753 (
            .O(N__31047),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    CascadeMux I__5752 (
            .O(N__31044),
            .I(N__31041));
    InMux I__5751 (
            .O(N__31041),
            .I(N__31035));
    InMux I__5750 (
            .O(N__31040),
            .I(N__31035));
    LocalMux I__5749 (
            .O(N__31035),
            .I(N__31031));
    InMux I__5748 (
            .O(N__31034),
            .I(N__31028));
    Span4Mux_v I__5747 (
            .O(N__31031),
            .I(N__31025));
    LocalMux I__5746 (
            .O(N__31028),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__5745 (
            .O(N__31025),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__5744 (
            .O(N__31020),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__5743 (
            .O(N__31017),
            .I(N__31011));
    InMux I__5742 (
            .O(N__31016),
            .I(N__31011));
    LocalMux I__5741 (
            .O(N__31011),
            .I(N__31007));
    InMux I__5740 (
            .O(N__31010),
            .I(N__31004));
    Span4Mux_h I__5739 (
            .O(N__31007),
            .I(N__31001));
    LocalMux I__5738 (
            .O(N__31004),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__5737 (
            .O(N__31001),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__5736 (
            .O(N__30996),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    CascadeMux I__5735 (
            .O(N__30993),
            .I(N__30990));
    InMux I__5734 (
            .O(N__30990),
            .I(N__30984));
    InMux I__5733 (
            .O(N__30989),
            .I(N__30984));
    LocalMux I__5732 (
            .O(N__30984),
            .I(N__30980));
    InMux I__5731 (
            .O(N__30983),
            .I(N__30977));
    Span4Mux_v I__5730 (
            .O(N__30980),
            .I(N__30974));
    LocalMux I__5729 (
            .O(N__30977),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__5728 (
            .O(N__30974),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__5727 (
            .O(N__30969),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__5726 (
            .O(N__30966),
            .I(N__30962));
    InMux I__5725 (
            .O(N__30965),
            .I(N__30959));
    LocalMux I__5724 (
            .O(N__30962),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__5723 (
            .O(N__30959),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__5722 (
            .O(N__30954),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__5721 (
            .O(N__30951),
            .I(N__30947));
    InMux I__5720 (
            .O(N__30950),
            .I(N__30944));
    LocalMux I__5719 (
            .O(N__30947),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__5718 (
            .O(N__30944),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__5717 (
            .O(N__30939),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__5716 (
            .O(N__30936),
            .I(N__30932));
    InMux I__5715 (
            .O(N__30935),
            .I(N__30929));
    LocalMux I__5714 (
            .O(N__30932),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__5713 (
            .O(N__30929),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__5712 (
            .O(N__30924),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__5711 (
            .O(N__30921),
            .I(N__30917));
    InMux I__5710 (
            .O(N__30920),
            .I(N__30914));
    LocalMux I__5709 (
            .O(N__30917),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__5708 (
            .O(N__30914),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__5707 (
            .O(N__30909),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__5706 (
            .O(N__30906),
            .I(N__30902));
    InMux I__5705 (
            .O(N__30905),
            .I(N__30899));
    LocalMux I__5704 (
            .O(N__30902),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__5703 (
            .O(N__30899),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__5702 (
            .O(N__30894),
            .I(bfn_12_11_0_));
    InMux I__5701 (
            .O(N__30891),
            .I(N__30887));
    InMux I__5700 (
            .O(N__30890),
            .I(N__30884));
    LocalMux I__5699 (
            .O(N__30887),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__5698 (
            .O(N__30884),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__5697 (
            .O(N__30879),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__5696 (
            .O(N__30876),
            .I(N__30872));
    InMux I__5695 (
            .O(N__30875),
            .I(N__30869));
    LocalMux I__5694 (
            .O(N__30872),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__5693 (
            .O(N__30869),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__5692 (
            .O(N__30864),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__5691 (
            .O(N__30861),
            .I(N__30857));
    InMux I__5690 (
            .O(N__30860),
            .I(N__30854));
    LocalMux I__5689 (
            .O(N__30857),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__5688 (
            .O(N__30854),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__5687 (
            .O(N__30849),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__5686 (
            .O(N__30846),
            .I(N__30843));
    LocalMux I__5685 (
            .O(N__30843),
            .I(N__30840));
    Span4Mux_h I__5684 (
            .O(N__30840),
            .I(N__30837));
    Odrv4 I__5683 (
            .O(N__30837),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ));
    CascadeMux I__5682 (
            .O(N__30834),
            .I(N__30831));
    InMux I__5681 (
            .O(N__30831),
            .I(N__30828));
    LocalMux I__5680 (
            .O(N__30828),
            .I(N__30825));
    Span4Mux_v I__5679 (
            .O(N__30825),
            .I(N__30822));
    Odrv4 I__5678 (
            .O(N__30822),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt26 ));
    InMux I__5677 (
            .O(N__30819),
            .I(N__30816));
    LocalMux I__5676 (
            .O(N__30816),
            .I(N__30813));
    Span4Mux_h I__5675 (
            .O(N__30813),
            .I(N__30810));
    Odrv4 I__5674 (
            .O(N__30810),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ));
    CascadeMux I__5673 (
            .O(N__30807),
            .I(N__30804));
    InMux I__5672 (
            .O(N__30804),
            .I(N__30801));
    LocalMux I__5671 (
            .O(N__30801),
            .I(N__30798));
    Span4Mux_v I__5670 (
            .O(N__30798),
            .I(N__30795));
    Odrv4 I__5669 (
            .O(N__30795),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt28 ));
    InMux I__5668 (
            .O(N__30792),
            .I(N__30789));
    LocalMux I__5667 (
            .O(N__30789),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    CascadeMux I__5666 (
            .O(N__30786),
            .I(N__30783));
    InMux I__5665 (
            .O(N__30783),
            .I(N__30779));
    InMux I__5664 (
            .O(N__30782),
            .I(N__30776));
    LocalMux I__5663 (
            .O(N__30779),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    LocalMux I__5662 (
            .O(N__30776),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    InMux I__5661 (
            .O(N__30771),
            .I(N__30768));
    LocalMux I__5660 (
            .O(N__30768),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__5659 (
            .O(N__30765),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ));
    InMux I__5658 (
            .O(N__30762),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    InMux I__5657 (
            .O(N__30759),
            .I(N__30753));
    InMux I__5656 (
            .O(N__30758),
            .I(N__30753));
    LocalMux I__5655 (
            .O(N__30753),
            .I(N__30750));
    Odrv12 I__5654 (
            .O(N__30750),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__5653 (
            .O(N__30747),
            .I(N__30744));
    LocalMux I__5652 (
            .O(N__30744),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    CascadeMux I__5651 (
            .O(N__30741),
            .I(N__30737));
    InMux I__5650 (
            .O(N__30740),
            .I(N__30733));
    InMux I__5649 (
            .O(N__30737),
            .I(N__30730));
    InMux I__5648 (
            .O(N__30736),
            .I(N__30727));
    LocalMux I__5647 (
            .O(N__30733),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__5646 (
            .O(N__30730),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__5645 (
            .O(N__30727),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__5644 (
            .O(N__30720),
            .I(N__30716));
    InMux I__5643 (
            .O(N__30719),
            .I(N__30713));
    LocalMux I__5642 (
            .O(N__30716),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__5641 (
            .O(N__30713),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__5640 (
            .O(N__30708),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__5639 (
            .O(N__30705),
            .I(N__30702));
    InMux I__5638 (
            .O(N__30702),
            .I(N__30699));
    LocalMux I__5637 (
            .O(N__30699),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ));
    InMux I__5636 (
            .O(N__30696),
            .I(N__30692));
    InMux I__5635 (
            .O(N__30695),
            .I(N__30689));
    LocalMux I__5634 (
            .O(N__30692),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__5633 (
            .O(N__30689),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__5632 (
            .O(N__30684),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__5631 (
            .O(N__30681),
            .I(N__30677));
    InMux I__5630 (
            .O(N__30680),
            .I(N__30674));
    LocalMux I__5629 (
            .O(N__30677),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__5628 (
            .O(N__30674),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__5627 (
            .O(N__30669),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__5626 (
            .O(N__30666),
            .I(N__30662));
    InMux I__5625 (
            .O(N__30665),
            .I(N__30659));
    LocalMux I__5624 (
            .O(N__30662),
            .I(N__30656));
    LocalMux I__5623 (
            .O(N__30659),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__5622 (
            .O(N__30656),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__5621 (
            .O(N__30651),
            .I(N__30648));
    LocalMux I__5620 (
            .O(N__30648),
            .I(N__30645));
    Span4Mux_h I__5619 (
            .O(N__30645),
            .I(N__30642));
    Span4Mux_h I__5618 (
            .O(N__30642),
            .I(N__30639));
    Odrv4 I__5617 (
            .O(N__30639),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__5616 (
            .O(N__30636),
            .I(N__30633));
    InMux I__5615 (
            .O(N__30633),
            .I(N__30630));
    LocalMux I__5614 (
            .O(N__30630),
            .I(N__30627));
    Odrv4 I__5613 (
            .O(N__30627),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__5612 (
            .O(N__30624),
            .I(N__30621));
    LocalMux I__5611 (
            .O(N__30621),
            .I(N__30617));
    InMux I__5610 (
            .O(N__30620),
            .I(N__30614));
    Span4Mux_v I__5609 (
            .O(N__30617),
            .I(N__30611));
    LocalMux I__5608 (
            .O(N__30614),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__5607 (
            .O(N__30611),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__5606 (
            .O(N__30606),
            .I(N__30603));
    InMux I__5605 (
            .O(N__30603),
            .I(N__30600));
    LocalMux I__5604 (
            .O(N__30600),
            .I(N__30597));
    Odrv12 I__5603 (
            .O(N__30597),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__5602 (
            .O(N__30594),
            .I(N__30591));
    LocalMux I__5601 (
            .O(N__30591),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__5600 (
            .O(N__30588),
            .I(N__30585));
    LocalMux I__5599 (
            .O(N__30585),
            .I(N__30582));
    Odrv12 I__5598 (
            .O(N__30582),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__5597 (
            .O(N__30579),
            .I(N__30575));
    InMux I__5596 (
            .O(N__30578),
            .I(N__30572));
    LocalMux I__5595 (
            .O(N__30575),
            .I(N__30569));
    LocalMux I__5594 (
            .O(N__30572),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__5593 (
            .O(N__30569),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__5592 (
            .O(N__30564),
            .I(N__30561));
    InMux I__5591 (
            .O(N__30561),
            .I(N__30558));
    LocalMux I__5590 (
            .O(N__30558),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__5589 (
            .O(N__30555),
            .I(N__30552));
    LocalMux I__5588 (
            .O(N__30552),
            .I(N__30549));
    Odrv4 I__5587 (
            .O(N__30549),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    CascadeMux I__5586 (
            .O(N__30546),
            .I(N__30543));
    InMux I__5585 (
            .O(N__30543),
            .I(N__30540));
    LocalMux I__5584 (
            .O(N__30540),
            .I(N__30537));
    Span4Mux_h I__5583 (
            .O(N__30537),
            .I(N__30534));
    Odrv4 I__5582 (
            .O(N__30534),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    InMux I__5581 (
            .O(N__30531),
            .I(N__30528));
    LocalMux I__5580 (
            .O(N__30528),
            .I(N__30525));
    Span4Mux_h I__5579 (
            .O(N__30525),
            .I(N__30522));
    Odrv4 I__5578 (
            .O(N__30522),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    CascadeMux I__5577 (
            .O(N__30519),
            .I(N__30516));
    InMux I__5576 (
            .O(N__30516),
            .I(N__30513));
    LocalMux I__5575 (
            .O(N__30513),
            .I(N__30510));
    Span4Mux_v I__5574 (
            .O(N__30510),
            .I(N__30507));
    Odrv4 I__5573 (
            .O(N__30507),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    InMux I__5572 (
            .O(N__30504),
            .I(N__30501));
    LocalMux I__5571 (
            .O(N__30501),
            .I(N__30498));
    Odrv4 I__5570 (
            .O(N__30498),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt20 ));
    CascadeMux I__5569 (
            .O(N__30495),
            .I(N__30492));
    InMux I__5568 (
            .O(N__30492),
            .I(N__30489));
    LocalMux I__5567 (
            .O(N__30489),
            .I(N__30486));
    Odrv4 I__5566 (
            .O(N__30486),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ));
    InMux I__5565 (
            .O(N__30483),
            .I(N__30480));
    LocalMux I__5564 (
            .O(N__30480),
            .I(N__30477));
    Span4Mux_h I__5563 (
            .O(N__30477),
            .I(N__30474));
    Odrv4 I__5562 (
            .O(N__30474),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ));
    CascadeMux I__5561 (
            .O(N__30471),
            .I(N__30468));
    InMux I__5560 (
            .O(N__30468),
            .I(N__30465));
    LocalMux I__5559 (
            .O(N__30465),
            .I(N__30462));
    Span4Mux_v I__5558 (
            .O(N__30462),
            .I(N__30459));
    Odrv4 I__5557 (
            .O(N__30459),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt22 ));
    InMux I__5556 (
            .O(N__30456),
            .I(N__30453));
    LocalMux I__5555 (
            .O(N__30453),
            .I(N__30450));
    Span4Mux_v I__5554 (
            .O(N__30450),
            .I(N__30447));
    Odrv4 I__5553 (
            .O(N__30447),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt24 ));
    CascadeMux I__5552 (
            .O(N__30444),
            .I(N__30441));
    InMux I__5551 (
            .O(N__30441),
            .I(N__30438));
    LocalMux I__5550 (
            .O(N__30438),
            .I(N__30435));
    Span4Mux_v I__5549 (
            .O(N__30435),
            .I(N__30432));
    Odrv4 I__5548 (
            .O(N__30432),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ));
    InMux I__5547 (
            .O(N__30429),
            .I(N__30425));
    InMux I__5546 (
            .O(N__30428),
            .I(N__30422));
    LocalMux I__5545 (
            .O(N__30425),
            .I(N__30419));
    LocalMux I__5544 (
            .O(N__30422),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__5543 (
            .O(N__30419),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__5542 (
            .O(N__30414),
            .I(N__30411));
    LocalMux I__5541 (
            .O(N__30411),
            .I(N__30408));
    Span4Mux_h I__5540 (
            .O(N__30408),
            .I(N__30405));
    Odrv4 I__5539 (
            .O(N__30405),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__5538 (
            .O(N__30402),
            .I(N__30399));
    InMux I__5537 (
            .O(N__30399),
            .I(N__30396));
    LocalMux I__5536 (
            .O(N__30396),
            .I(N__30393));
    Odrv4 I__5535 (
            .O(N__30393),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__5534 (
            .O(N__30390),
            .I(N__30387));
    LocalMux I__5533 (
            .O(N__30387),
            .I(N__30384));
    Odrv12 I__5532 (
            .O(N__30384),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__5531 (
            .O(N__30381),
            .I(N__30377));
    InMux I__5530 (
            .O(N__30380),
            .I(N__30374));
    LocalMux I__5529 (
            .O(N__30377),
            .I(N__30371));
    LocalMux I__5528 (
            .O(N__30374),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__5527 (
            .O(N__30371),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__5526 (
            .O(N__30366),
            .I(N__30363));
    InMux I__5525 (
            .O(N__30363),
            .I(N__30360));
    LocalMux I__5524 (
            .O(N__30360),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__5523 (
            .O(N__30357),
            .I(N__30353));
    InMux I__5522 (
            .O(N__30356),
            .I(N__30350));
    LocalMux I__5521 (
            .O(N__30353),
            .I(N__30347));
    LocalMux I__5520 (
            .O(N__30350),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__5519 (
            .O(N__30347),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__5518 (
            .O(N__30342),
            .I(N__30339));
    LocalMux I__5517 (
            .O(N__30339),
            .I(N__30336));
    Span4Mux_v I__5516 (
            .O(N__30336),
            .I(N__30333));
    Span4Mux_v I__5515 (
            .O(N__30333),
            .I(N__30330));
    Span4Mux_h I__5514 (
            .O(N__30330),
            .I(N__30327));
    Odrv4 I__5513 (
            .O(N__30327),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__5512 (
            .O(N__30324),
            .I(N__30321));
    InMux I__5511 (
            .O(N__30321),
            .I(N__30318));
    LocalMux I__5510 (
            .O(N__30318),
            .I(N__30315));
    Odrv4 I__5509 (
            .O(N__30315),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__5508 (
            .O(N__30312),
            .I(N__30309));
    LocalMux I__5507 (
            .O(N__30309),
            .I(N__30306));
    Span4Mux_h I__5506 (
            .O(N__30306),
            .I(N__30303));
    Odrv4 I__5505 (
            .O(N__30303),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__5504 (
            .O(N__30300),
            .I(N__30297));
    LocalMux I__5503 (
            .O(N__30297),
            .I(N__30293));
    InMux I__5502 (
            .O(N__30296),
            .I(N__30290));
    Span4Mux_v I__5501 (
            .O(N__30293),
            .I(N__30287));
    LocalMux I__5500 (
            .O(N__30290),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__5499 (
            .O(N__30287),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__5498 (
            .O(N__30282),
            .I(N__30279));
    InMux I__5497 (
            .O(N__30279),
            .I(N__30276));
    LocalMux I__5496 (
            .O(N__30276),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__5495 (
            .O(N__30273),
            .I(N__30270));
    LocalMux I__5494 (
            .O(N__30270),
            .I(N__30267));
    Span4Mux_v I__5493 (
            .O(N__30267),
            .I(N__30264));
    Odrv4 I__5492 (
            .O(N__30264),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__5491 (
            .O(N__30261),
            .I(N__30257));
    InMux I__5490 (
            .O(N__30260),
            .I(N__30254));
    LocalMux I__5489 (
            .O(N__30257),
            .I(N__30251));
    LocalMux I__5488 (
            .O(N__30254),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__5487 (
            .O(N__30251),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__5486 (
            .O(N__30246),
            .I(N__30243));
    InMux I__5485 (
            .O(N__30243),
            .I(N__30240));
    LocalMux I__5484 (
            .O(N__30240),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__5483 (
            .O(N__30237),
            .I(N__30234));
    LocalMux I__5482 (
            .O(N__30234),
            .I(N__30231));
    Span4Mux_h I__5481 (
            .O(N__30231),
            .I(N__30228));
    Odrv4 I__5480 (
            .O(N__30228),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__5479 (
            .O(N__30225),
            .I(N__30222));
    LocalMux I__5478 (
            .O(N__30222),
            .I(N__30218));
    InMux I__5477 (
            .O(N__30221),
            .I(N__30215));
    Span4Mux_v I__5476 (
            .O(N__30218),
            .I(N__30212));
    LocalMux I__5475 (
            .O(N__30215),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__5474 (
            .O(N__30212),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__5473 (
            .O(N__30207),
            .I(N__30204));
    InMux I__5472 (
            .O(N__30204),
            .I(N__30201));
    LocalMux I__5471 (
            .O(N__30201),
            .I(N__30198));
    Odrv4 I__5470 (
            .O(N__30198),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__5469 (
            .O(N__30195),
            .I(N__30192));
    LocalMux I__5468 (
            .O(N__30192),
            .I(N__30189));
    Odrv12 I__5467 (
            .O(N__30189),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__5466 (
            .O(N__30186),
            .I(N__30182));
    InMux I__5465 (
            .O(N__30185),
            .I(N__30179));
    LocalMux I__5464 (
            .O(N__30182),
            .I(N__30176));
    LocalMux I__5463 (
            .O(N__30179),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__5462 (
            .O(N__30176),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__5461 (
            .O(N__30171),
            .I(N__30168));
    InMux I__5460 (
            .O(N__30168),
            .I(N__30165));
    LocalMux I__5459 (
            .O(N__30165),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__5458 (
            .O(N__30162),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ));
    InMux I__5457 (
            .O(N__30159),
            .I(N__30156));
    LocalMux I__5456 (
            .O(N__30156),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ));
    InMux I__5455 (
            .O(N__30153),
            .I(N__30141));
    InMux I__5454 (
            .O(N__30152),
            .I(N__30141));
    InMux I__5453 (
            .O(N__30151),
            .I(N__30141));
    InMux I__5452 (
            .O(N__30150),
            .I(N__30141));
    LocalMux I__5451 (
            .O(N__30141),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    CascadeMux I__5450 (
            .O(N__30138),
            .I(N__30133));
    CascadeMux I__5449 (
            .O(N__30137),
            .I(N__30130));
    InMux I__5448 (
            .O(N__30136),
            .I(N__30125));
    InMux I__5447 (
            .O(N__30133),
            .I(N__30116));
    InMux I__5446 (
            .O(N__30130),
            .I(N__30116));
    InMux I__5445 (
            .O(N__30129),
            .I(N__30116));
    InMux I__5444 (
            .O(N__30128),
            .I(N__30116));
    LocalMux I__5443 (
            .O(N__30125),
            .I(N__30113));
    LocalMux I__5442 (
            .O(N__30116),
            .I(N__30108));
    Span4Mux_v I__5441 (
            .O(N__30113),
            .I(N__30108));
    Odrv4 I__5440 (
            .O(N__30108),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__5439 (
            .O(N__30105),
            .I(N__30102));
    LocalMux I__5438 (
            .O(N__30102),
            .I(N__30099));
    Span4Mux_h I__5437 (
            .O(N__30099),
            .I(N__30096));
    Odrv4 I__5436 (
            .O(N__30096),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__5435 (
            .O(N__30093),
            .I(N__30090));
    InMux I__5434 (
            .O(N__30090),
            .I(N__30087));
    LocalMux I__5433 (
            .O(N__30087),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__5432 (
            .O(N__30084),
            .I(N__30081));
    LocalMux I__5431 (
            .O(N__30081),
            .I(N__30078));
    Span4Mux_h I__5430 (
            .O(N__30078),
            .I(N__30075));
    Odrv4 I__5429 (
            .O(N__30075),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__5428 (
            .O(N__30072),
            .I(N__30068));
    InMux I__5427 (
            .O(N__30071),
            .I(N__30065));
    LocalMux I__5426 (
            .O(N__30068),
            .I(N__30062));
    LocalMux I__5425 (
            .O(N__30065),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__5424 (
            .O(N__30062),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__5423 (
            .O(N__30057),
            .I(N__30054));
    InMux I__5422 (
            .O(N__30054),
            .I(N__30051));
    LocalMux I__5421 (
            .O(N__30051),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__5420 (
            .O(N__30048),
            .I(N__30045));
    LocalMux I__5419 (
            .O(N__30045),
            .I(N__30042));
    Span4Mux_h I__5418 (
            .O(N__30042),
            .I(N__30039));
    Odrv4 I__5417 (
            .O(N__30039),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__5416 (
            .O(N__30036),
            .I(N__30032));
    CascadeMux I__5415 (
            .O(N__30035),
            .I(N__30029));
    LocalMux I__5414 (
            .O(N__30032),
            .I(N__30026));
    InMux I__5413 (
            .O(N__30029),
            .I(N__30023));
    Span4Mux_v I__5412 (
            .O(N__30026),
            .I(N__30020));
    LocalMux I__5411 (
            .O(N__30023),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__5410 (
            .O(N__30020),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__5409 (
            .O(N__30015),
            .I(N__30012));
    InMux I__5408 (
            .O(N__30012),
            .I(N__30009));
    LocalMux I__5407 (
            .O(N__30009),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__5406 (
            .O(N__30006),
            .I(N__30003));
    LocalMux I__5405 (
            .O(N__30003),
            .I(N__30000));
    Span4Mux_v I__5404 (
            .O(N__30000),
            .I(N__29997));
    Odrv4 I__5403 (
            .O(N__29997),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__5402 (
            .O(N__29994),
            .I(N__29990));
    InMux I__5401 (
            .O(N__29993),
            .I(N__29987));
    LocalMux I__5400 (
            .O(N__29990),
            .I(N__29984));
    LocalMux I__5399 (
            .O(N__29987),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__5398 (
            .O(N__29984),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__5397 (
            .O(N__29979),
            .I(N__29976));
    InMux I__5396 (
            .O(N__29976),
            .I(N__29973));
    LocalMux I__5395 (
            .O(N__29973),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__5394 (
            .O(N__29970),
            .I(N__29966));
    InMux I__5393 (
            .O(N__29969),
            .I(N__29963));
    LocalMux I__5392 (
            .O(N__29966),
            .I(N__29960));
    LocalMux I__5391 (
            .O(N__29963),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__5390 (
            .O(N__29960),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__5389 (
            .O(N__29955),
            .I(N__29952));
    LocalMux I__5388 (
            .O(N__29952),
            .I(N__29949));
    Odrv4 I__5387 (
            .O(N__29949),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__5386 (
            .O(N__29946),
            .I(N__29943));
    InMux I__5385 (
            .O(N__29943),
            .I(N__29940));
    LocalMux I__5384 (
            .O(N__29940),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__5383 (
            .O(N__29937),
            .I(N__29933));
    InMux I__5382 (
            .O(N__29936),
            .I(N__29929));
    LocalMux I__5381 (
            .O(N__29933),
            .I(N__29926));
    InMux I__5380 (
            .O(N__29932),
            .I(N__29923));
    LocalMux I__5379 (
            .O(N__29929),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv4 I__5378 (
            .O(N__29926),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__5377 (
            .O(N__29923),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    CascadeMux I__5376 (
            .O(N__29916),
            .I(N__29913));
    InMux I__5375 (
            .O(N__29913),
            .I(N__29910));
    LocalMux I__5374 (
            .O(N__29910),
            .I(N__29907));
    Span4Mux_h I__5373 (
            .O(N__29907),
            .I(N__29903));
    InMux I__5372 (
            .O(N__29906),
            .I(N__29900));
    Odrv4 I__5371 (
            .O(N__29903),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    LocalMux I__5370 (
            .O(N__29900),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__5369 (
            .O(N__29895),
            .I(N__29892));
    LocalMux I__5368 (
            .O(N__29892),
            .I(N__29889));
    Odrv12 I__5367 (
            .O(N__29889),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    CascadeMux I__5366 (
            .O(N__29886),
            .I(N__29882));
    InMux I__5365 (
            .O(N__29885),
            .I(N__29877));
    InMux I__5364 (
            .O(N__29882),
            .I(N__29874));
    CascadeMux I__5363 (
            .O(N__29881),
            .I(N__29869));
    CascadeMux I__5362 (
            .O(N__29880),
            .I(N__29863));
    LocalMux I__5361 (
            .O(N__29877),
            .I(N__29858));
    LocalMux I__5360 (
            .O(N__29874),
            .I(N__29858));
    InMux I__5359 (
            .O(N__29873),
            .I(N__29855));
    CascadeMux I__5358 (
            .O(N__29872),
            .I(N__29852));
    InMux I__5357 (
            .O(N__29869),
            .I(N__29843));
    InMux I__5356 (
            .O(N__29868),
            .I(N__29843));
    InMux I__5355 (
            .O(N__29867),
            .I(N__29843));
    InMux I__5354 (
            .O(N__29866),
            .I(N__29843));
    InMux I__5353 (
            .O(N__29863),
            .I(N__29840));
    Span4Mux_h I__5352 (
            .O(N__29858),
            .I(N__29835));
    LocalMux I__5351 (
            .O(N__29855),
            .I(N__29835));
    InMux I__5350 (
            .O(N__29852),
            .I(N__29832));
    LocalMux I__5349 (
            .O(N__29843),
            .I(N__29824));
    LocalMux I__5348 (
            .O(N__29840),
            .I(N__29824));
    Span4Mux_v I__5347 (
            .O(N__29835),
            .I(N__29821));
    LocalMux I__5346 (
            .O(N__29832),
            .I(N__29818));
    InMux I__5345 (
            .O(N__29831),
            .I(N__29815));
    InMux I__5344 (
            .O(N__29830),
            .I(N__29810));
    InMux I__5343 (
            .O(N__29829),
            .I(N__29810));
    Span4Mux_v I__5342 (
            .O(N__29824),
            .I(N__29807));
    Span4Mux_s2_v I__5341 (
            .O(N__29821),
            .I(N__29804));
    Odrv4 I__5340 (
            .O(N__29818),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    LocalMux I__5339 (
            .O(N__29815),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    LocalMux I__5338 (
            .O(N__29810),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__5337 (
            .O(N__29807),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__5336 (
            .O(N__29804),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    InMux I__5335 (
            .O(N__29793),
            .I(N__29790));
    LocalMux I__5334 (
            .O(N__29790),
            .I(N__29787));
    Odrv12 I__5333 (
            .O(N__29787),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    CascadeMux I__5332 (
            .O(N__29784),
            .I(N__29781));
    InMux I__5331 (
            .O(N__29781),
            .I(N__29777));
    InMux I__5330 (
            .O(N__29780),
            .I(N__29773));
    LocalMux I__5329 (
            .O(N__29777),
            .I(N__29770));
    InMux I__5328 (
            .O(N__29776),
            .I(N__29767));
    LocalMux I__5327 (
            .O(N__29773),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    Odrv4 I__5326 (
            .O(N__29770),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__5325 (
            .O(N__29767),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    InMux I__5324 (
            .O(N__29760),
            .I(N__29757));
    LocalMux I__5323 (
            .O(N__29757),
            .I(N__29754));
    Span4Mux_v I__5322 (
            .O(N__29754),
            .I(N__29750));
    InMux I__5321 (
            .O(N__29753),
            .I(N__29747));
    Odrv4 I__5320 (
            .O(N__29750),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    LocalMux I__5319 (
            .O(N__29747),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    InMux I__5318 (
            .O(N__29742),
            .I(N__29739));
    LocalMux I__5317 (
            .O(N__29739),
            .I(N__29736));
    Odrv12 I__5316 (
            .O(N__29736),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    InMux I__5315 (
            .O(N__29733),
            .I(N__29729));
    InMux I__5314 (
            .O(N__29732),
            .I(N__29726));
    LocalMux I__5313 (
            .O(N__29729),
            .I(N__29723));
    LocalMux I__5312 (
            .O(N__29726),
            .I(N__29720));
    Span4Mux_h I__5311 (
            .O(N__29723),
            .I(N__29715));
    Span4Mux_h I__5310 (
            .O(N__29720),
            .I(N__29715));
    Span4Mux_v I__5309 (
            .O(N__29715),
            .I(N__29710));
    InMux I__5308 (
            .O(N__29714),
            .I(N__29707));
    InMux I__5307 (
            .O(N__29713),
            .I(N__29704));
    Span4Mux_v I__5306 (
            .O(N__29710),
            .I(N__29701));
    LocalMux I__5305 (
            .O(N__29707),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__5304 (
            .O(N__29704),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__5303 (
            .O(N__29701),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    ClkMux I__5302 (
            .O(N__29694),
            .I(N__29688));
    ClkMux I__5301 (
            .O(N__29693),
            .I(N__29688));
    GlobalMux I__5300 (
            .O(N__29688),
            .I(N__29685));
    gio2CtrlBuf I__5299 (
            .O(N__29685),
            .I(delay_hc_input_c_g));
    InMux I__5298 (
            .O(N__29682),
            .I(N__29677));
    InMux I__5297 (
            .O(N__29681),
            .I(N__29673));
    CascadeMux I__5296 (
            .O(N__29680),
            .I(N__29670));
    LocalMux I__5295 (
            .O(N__29677),
            .I(N__29667));
    InMux I__5294 (
            .O(N__29676),
            .I(N__29664));
    LocalMux I__5293 (
            .O(N__29673),
            .I(N__29661));
    InMux I__5292 (
            .O(N__29670),
            .I(N__29658));
    Span4Mux_v I__5291 (
            .O(N__29667),
            .I(N__29655));
    LocalMux I__5290 (
            .O(N__29664),
            .I(N__29648));
    Span4Mux_v I__5289 (
            .O(N__29661),
            .I(N__29648));
    LocalMux I__5288 (
            .O(N__29658),
            .I(N__29648));
    Span4Mux_h I__5287 (
            .O(N__29655),
            .I(N__29645));
    Span4Mux_v I__5286 (
            .O(N__29648),
            .I(N__29642));
    Odrv4 I__5285 (
            .O(N__29645),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__5284 (
            .O(N__29642),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__5283 (
            .O(N__29637),
            .I(N__29632));
    InMux I__5282 (
            .O(N__29636),
            .I(N__29629));
    InMux I__5281 (
            .O(N__29635),
            .I(N__29626));
    LocalMux I__5280 (
            .O(N__29632),
            .I(N__29623));
    LocalMux I__5279 (
            .O(N__29629),
            .I(N__29620));
    LocalMux I__5278 (
            .O(N__29626),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    Odrv12 I__5277 (
            .O(N__29623),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    Odrv4 I__5276 (
            .O(N__29620),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    InMux I__5275 (
            .O(N__29613),
            .I(N__29610));
    LocalMux I__5274 (
            .O(N__29610),
            .I(N__29607));
    Span4Mux_h I__5273 (
            .O(N__29607),
            .I(N__29604));
    Span4Mux_v I__5272 (
            .O(N__29604),
            .I(N__29601));
    Odrv4 I__5271 (
            .O(N__29601),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    CascadeMux I__5270 (
            .O(N__29598),
            .I(N__29595));
    InMux I__5269 (
            .O(N__29595),
            .I(N__29592));
    LocalMux I__5268 (
            .O(N__29592),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    InMux I__5267 (
            .O(N__29589),
            .I(N__29583));
    InMux I__5266 (
            .O(N__29588),
            .I(N__29583));
    LocalMux I__5265 (
            .O(N__29583),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    InMux I__5264 (
            .O(N__29580),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__5263 (
            .O(N__29577),
            .I(N__29574));
    LocalMux I__5262 (
            .O(N__29574),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__5261 (
            .O(N__29571),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__5260 (
            .O(N__29568),
            .I(N__29565));
    LocalMux I__5259 (
            .O(N__29565),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    InMux I__5258 (
            .O(N__29562),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    InMux I__5257 (
            .O(N__29559),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__5256 (
            .O(N__29556),
            .I(N__29553));
    LocalMux I__5255 (
            .O(N__29553),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__5254 (
            .O(N__29550),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__5253 (
            .O(N__29547),
            .I(N__29544));
    LocalMux I__5252 (
            .O(N__29544),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    InMux I__5251 (
            .O(N__29541),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    InMux I__5250 (
            .O(N__29538),
            .I(N__29535));
    LocalMux I__5249 (
            .O(N__29535),
            .I(N__29532));
    Span4Mux_h I__5248 (
            .O(N__29532),
            .I(N__29529));
    Odrv4 I__5247 (
            .O(N__29529),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__5246 (
            .O(N__29526),
            .I(bfn_11_25_0_));
    InMux I__5245 (
            .O(N__29523),
            .I(N__29520));
    LocalMux I__5244 (
            .O(N__29520),
            .I(N__29517));
    Span4Mux_h I__5243 (
            .O(N__29517),
            .I(N__29514));
    Odrv4 I__5242 (
            .O(N__29514),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    InMux I__5241 (
            .O(N__29511),
            .I(N__29508));
    LocalMux I__5240 (
            .O(N__29508),
            .I(N__29505));
    Span4Mux_h I__5239 (
            .O(N__29505),
            .I(N__29502));
    Odrv4 I__5238 (
            .O(N__29502),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ));
    InMux I__5237 (
            .O(N__29499),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    InMux I__5236 (
            .O(N__29496),
            .I(N__29493));
    LocalMux I__5235 (
            .O(N__29493),
            .I(N__29490));
    Odrv12 I__5234 (
            .O(N__29490),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    InMux I__5233 (
            .O(N__29487),
            .I(N__29484));
    LocalMux I__5232 (
            .O(N__29484),
            .I(N__29481));
    Odrv12 I__5231 (
            .O(N__29481),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__5230 (
            .O(N__29478),
            .I(N__29475));
    LocalMux I__5229 (
            .O(N__29475),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__5228 (
            .O(N__29472),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__5227 (
            .O(N__29469),
            .I(N__29466));
    LocalMux I__5226 (
            .O(N__29466),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__5225 (
            .O(N__29463),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__5224 (
            .O(N__29460),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__5223 (
            .O(N__29457),
            .I(N__29454));
    LocalMux I__5222 (
            .O(N__29454),
            .I(N__29451));
    Span12Mux_v I__5221 (
            .O(N__29451),
            .I(N__29448));
    Odrv12 I__5220 (
            .O(N__29448),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__5219 (
            .O(N__29445),
            .I(N__29442));
    LocalMux I__5218 (
            .O(N__29442),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__5217 (
            .O(N__29439),
            .I(N__29436));
    LocalMux I__5216 (
            .O(N__29436),
            .I(N__29433));
    Span4Mux_v I__5215 (
            .O(N__29433),
            .I(N__29430));
    Span4Mux_h I__5214 (
            .O(N__29430),
            .I(N__29427));
    Odrv4 I__5213 (
            .O(N__29427),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__5212 (
            .O(N__29424),
            .I(N__29421));
    LocalMux I__5211 (
            .O(N__29421),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__5210 (
            .O(N__29418),
            .I(N__29415));
    LocalMux I__5209 (
            .O(N__29415),
            .I(N__29412));
    Span4Mux_h I__5208 (
            .O(N__29412),
            .I(N__29409));
    Span4Mux_v I__5207 (
            .O(N__29409),
            .I(N__29406));
    Odrv4 I__5206 (
            .O(N__29406),
            .I(\current_shift_inst.control_input_axb_4 ));
    IoInMux I__5205 (
            .O(N__29403),
            .I(N__29400));
    LocalMux I__5204 (
            .O(N__29400),
            .I(N__29397));
    Span4Mux_s3_v I__5203 (
            .O(N__29397),
            .I(N__29394));
    Span4Mux_v I__5202 (
            .O(N__29394),
            .I(N__29391));
    Odrv4 I__5201 (
            .O(N__29391),
            .I(s3_phy_c));
    InMux I__5200 (
            .O(N__29388),
            .I(N__29385));
    LocalMux I__5199 (
            .O(N__29385),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    InMux I__5198 (
            .O(N__29382),
            .I(N__29379));
    LocalMux I__5197 (
            .O(N__29379),
            .I(N__29376));
    Span4Mux_h I__5196 (
            .O(N__29376),
            .I(N__29373));
    Odrv4 I__5195 (
            .O(N__29373),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__5194 (
            .O(N__29370),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    InMux I__5193 (
            .O(N__29367),
            .I(N__29364));
    LocalMux I__5192 (
            .O(N__29364),
            .I(N__29361));
    Span4Mux_v I__5191 (
            .O(N__29361),
            .I(N__29358));
    Odrv4 I__5190 (
            .O(N__29358),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__5189 (
            .O(N__29355),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__5188 (
            .O(N__29352),
            .I(N__29349));
    LocalMux I__5187 (
            .O(N__29349),
            .I(N__29346));
    Span4Mux_h I__5186 (
            .O(N__29346),
            .I(N__29343));
    Odrv4 I__5185 (
            .O(N__29343),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__5184 (
            .O(N__29340),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__5183 (
            .O(N__29337),
            .I(N__29334));
    LocalMux I__5182 (
            .O(N__29334),
            .I(N__29331));
    Span4Mux_h I__5181 (
            .O(N__29331),
            .I(N__29328));
    Odrv4 I__5180 (
            .O(N__29328),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__5179 (
            .O(N__29325),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__5178 (
            .O(N__29322),
            .I(bfn_11_20_0_));
    InMux I__5177 (
            .O(N__29319),
            .I(N__29316));
    LocalMux I__5176 (
            .O(N__29316),
            .I(N__29313));
    Span4Mux_h I__5175 (
            .O(N__29313),
            .I(N__29310));
    Odrv4 I__5174 (
            .O(N__29310),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__5173 (
            .O(N__29307),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__5172 (
            .O(N__29304),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__5171 (
            .O(N__29301),
            .I(N__29298));
    LocalMux I__5170 (
            .O(N__29298),
            .I(N__29295));
    Span4Mux_h I__5169 (
            .O(N__29295),
            .I(N__29292));
    Odrv4 I__5168 (
            .O(N__29292),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__5167 (
            .O(N__29289),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__5166 (
            .O(N__29286),
            .I(N__29283));
    LocalMux I__5165 (
            .O(N__29283),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__5164 (
            .O(N__29280),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    CascadeMux I__5163 (
            .O(N__29277),
            .I(N__29274));
    InMux I__5162 (
            .O(N__29274),
            .I(N__29271));
    LocalMux I__5161 (
            .O(N__29271),
            .I(N__29268));
    Odrv4 I__5160 (
            .O(N__29268),
            .I(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ));
    InMux I__5159 (
            .O(N__29265),
            .I(N__29262));
    LocalMux I__5158 (
            .O(N__29262),
            .I(N__29259));
    Odrv4 I__5157 (
            .O(N__29259),
            .I(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ));
    InMux I__5156 (
            .O(N__29256),
            .I(N__29253));
    LocalMux I__5155 (
            .O(N__29253),
            .I(N__29250));
    Span4Mux_v I__5154 (
            .O(N__29250),
            .I(N__29247));
    Odrv4 I__5153 (
            .O(N__29247),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__5152 (
            .O(N__29244),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    CascadeMux I__5151 (
            .O(N__29241),
            .I(N__29238));
    InMux I__5150 (
            .O(N__29238),
            .I(N__29235));
    LocalMux I__5149 (
            .O(N__29235),
            .I(N__29232));
    Odrv4 I__5148 (
            .O(N__29232),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    CascadeMux I__5147 (
            .O(N__29229),
            .I(N__29226));
    InMux I__5146 (
            .O(N__29226),
            .I(N__29223));
    LocalMux I__5145 (
            .O(N__29223),
            .I(N__29220));
    Odrv4 I__5144 (
            .O(N__29220),
            .I(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ));
    InMux I__5143 (
            .O(N__29217),
            .I(N__29214));
    LocalMux I__5142 (
            .O(N__29214),
            .I(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ));
    InMux I__5141 (
            .O(N__29211),
            .I(N__29208));
    LocalMux I__5140 (
            .O(N__29208),
            .I(N__29205));
    Odrv4 I__5139 (
            .O(N__29205),
            .I(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ));
    InMux I__5138 (
            .O(N__29202),
            .I(N__29198));
    InMux I__5137 (
            .O(N__29201),
            .I(N__29195));
    LocalMux I__5136 (
            .O(N__29198),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__5135 (
            .O(N__29195),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    CascadeMux I__5134 (
            .O(N__29190),
            .I(N__29187));
    InMux I__5133 (
            .O(N__29187),
            .I(N__29184));
    LocalMux I__5132 (
            .O(N__29184),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__5131 (
            .O(N__29181),
            .I(N__29178));
    LocalMux I__5130 (
            .O(N__29178),
            .I(N__29175));
    Span4Mux_v I__5129 (
            .O(N__29175),
            .I(N__29172));
    Odrv4 I__5128 (
            .O(N__29172),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    CascadeMux I__5127 (
            .O(N__29169),
            .I(N__29166));
    InMux I__5126 (
            .O(N__29166),
            .I(N__29163));
    LocalMux I__5125 (
            .O(N__29163),
            .I(N__29159));
    InMux I__5124 (
            .O(N__29162),
            .I(N__29156));
    Odrv12 I__5123 (
            .O(N__29159),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    LocalMux I__5122 (
            .O(N__29156),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    InMux I__5121 (
            .O(N__29151),
            .I(N__29148));
    LocalMux I__5120 (
            .O(N__29148),
            .I(N__29145));
    Odrv12 I__5119 (
            .O(N__29145),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__5118 (
            .O(N__29142),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ));
    InMux I__5117 (
            .O(N__29139),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    InMux I__5116 (
            .O(N__29136),
            .I(N__29133));
    LocalMux I__5115 (
            .O(N__29133),
            .I(N__29130));
    Sp12to4 I__5114 (
            .O(N__29130),
            .I(N__29127));
    Span12Mux_v I__5113 (
            .O(N__29127),
            .I(N__29124));
    Odrv12 I__5112 (
            .O(N__29124),
            .I(il_max_comp1_D1));
    InMux I__5111 (
            .O(N__29121),
            .I(N__29118));
    LocalMux I__5110 (
            .O(N__29118),
            .I(N__29115));
    Odrv4 I__5109 (
            .O(N__29115),
            .I(il_min_comp1_D1));
    CascadeMux I__5108 (
            .O(N__29112),
            .I(N__29109));
    InMux I__5107 (
            .O(N__29109),
            .I(N__29106));
    LocalMux I__5106 (
            .O(N__29106),
            .I(N__29103));
    Odrv12 I__5105 (
            .O(N__29103),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    InMux I__5104 (
            .O(N__29100),
            .I(N__29097));
    LocalMux I__5103 (
            .O(N__29097),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__5102 (
            .O(N__29094),
            .I(N__29091));
    LocalMux I__5101 (
            .O(N__29091),
            .I(N__29088));
    Sp12to4 I__5100 (
            .O(N__29088),
            .I(N__29085));
    Odrv12 I__5099 (
            .O(N__29085),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    CascadeMux I__5098 (
            .O(N__29082),
            .I(N__29079));
    InMux I__5097 (
            .O(N__29079),
            .I(N__29076));
    LocalMux I__5096 (
            .O(N__29076),
            .I(N__29073));
    Span4Mux_h I__5095 (
            .O(N__29073),
            .I(N__29070));
    Odrv4 I__5094 (
            .O(N__29070),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    InMux I__5093 (
            .O(N__29067),
            .I(N__29064));
    LocalMux I__5092 (
            .O(N__29064),
            .I(N__29061));
    Span4Mux_v I__5091 (
            .O(N__29061),
            .I(N__29058));
    Odrv4 I__5090 (
            .O(N__29058),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    CascadeMux I__5089 (
            .O(N__29055),
            .I(N__29052));
    InMux I__5088 (
            .O(N__29052),
            .I(N__29049));
    LocalMux I__5087 (
            .O(N__29049),
            .I(N__29046));
    Span4Mux_v I__5086 (
            .O(N__29046),
            .I(N__29043));
    Odrv4 I__5085 (
            .O(N__29043),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    InMux I__5084 (
            .O(N__29040),
            .I(N__29037));
    LocalMux I__5083 (
            .O(N__29037),
            .I(N__29034));
    Odrv4 I__5082 (
            .O(N__29034),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ));
    CascadeMux I__5081 (
            .O(N__29031),
            .I(N__29028));
    InMux I__5080 (
            .O(N__29028),
            .I(N__29025));
    LocalMux I__5079 (
            .O(N__29025),
            .I(N__29022));
    Odrv12 I__5078 (
            .O(N__29022),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt20 ));
    InMux I__5077 (
            .O(N__29019),
            .I(N__29016));
    LocalMux I__5076 (
            .O(N__29016),
            .I(N__29013));
    Odrv4 I__5075 (
            .O(N__29013),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ));
    CascadeMux I__5074 (
            .O(N__29010),
            .I(N__29007));
    InMux I__5073 (
            .O(N__29007),
            .I(N__29004));
    LocalMux I__5072 (
            .O(N__29004),
            .I(N__29001));
    Span4Mux_h I__5071 (
            .O(N__29001),
            .I(N__28998));
    Odrv4 I__5070 (
            .O(N__28998),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt22 ));
    InMux I__5069 (
            .O(N__28995),
            .I(N__28992));
    LocalMux I__5068 (
            .O(N__28992),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ));
    CascadeMux I__5067 (
            .O(N__28989),
            .I(N__28986));
    InMux I__5066 (
            .O(N__28986),
            .I(N__28983));
    LocalMux I__5065 (
            .O(N__28983),
            .I(N__28980));
    Odrv4 I__5064 (
            .O(N__28980),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt24 ));
    InMux I__5063 (
            .O(N__28977),
            .I(N__28974));
    LocalMux I__5062 (
            .O(N__28974),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ));
    CascadeMux I__5061 (
            .O(N__28971),
            .I(N__28968));
    InMux I__5060 (
            .O(N__28968),
            .I(N__28965));
    LocalMux I__5059 (
            .O(N__28965),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt26 ));
    InMux I__5058 (
            .O(N__28962),
            .I(N__28959));
    LocalMux I__5057 (
            .O(N__28959),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ));
    CascadeMux I__5056 (
            .O(N__28956),
            .I(N__28953));
    InMux I__5055 (
            .O(N__28953),
            .I(N__28950));
    LocalMux I__5054 (
            .O(N__28950),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt28 ));
    InMux I__5053 (
            .O(N__28947),
            .I(N__28944));
    LocalMux I__5052 (
            .O(N__28944),
            .I(N__28941));
    Odrv4 I__5051 (
            .O(N__28941),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__5050 (
            .O(N__28938),
            .I(N__28935));
    InMux I__5049 (
            .O(N__28935),
            .I(N__28932));
    LocalMux I__5048 (
            .O(N__28932),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__5047 (
            .O(N__28929),
            .I(N__28926));
    LocalMux I__5046 (
            .O(N__28926),
            .I(N__28923));
    Span4Mux_v I__5045 (
            .O(N__28923),
            .I(N__28920));
    Odrv4 I__5044 (
            .O(N__28920),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__5043 (
            .O(N__28917),
            .I(N__28914));
    InMux I__5042 (
            .O(N__28914),
            .I(N__28911));
    LocalMux I__5041 (
            .O(N__28911),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__5040 (
            .O(N__28908),
            .I(N__28905));
    LocalMux I__5039 (
            .O(N__28905),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__5038 (
            .O(N__28902),
            .I(N__28899));
    InMux I__5037 (
            .O(N__28899),
            .I(N__28896));
    LocalMux I__5036 (
            .O(N__28896),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__5035 (
            .O(N__28893),
            .I(N__28890));
    LocalMux I__5034 (
            .O(N__28890),
            .I(N__28887));
    Span4Mux_h I__5033 (
            .O(N__28887),
            .I(N__28884));
    Odrv4 I__5032 (
            .O(N__28884),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__5031 (
            .O(N__28881),
            .I(N__28878));
    InMux I__5030 (
            .O(N__28878),
            .I(N__28875));
    LocalMux I__5029 (
            .O(N__28875),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__5028 (
            .O(N__28872),
            .I(N__28869));
    LocalMux I__5027 (
            .O(N__28869),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__5026 (
            .O(N__28866),
            .I(N__28863));
    InMux I__5025 (
            .O(N__28863),
            .I(N__28860));
    LocalMux I__5024 (
            .O(N__28860),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__5023 (
            .O(N__28857),
            .I(N__28854));
    LocalMux I__5022 (
            .O(N__28854),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__5021 (
            .O(N__28851),
            .I(N__28848));
    InMux I__5020 (
            .O(N__28848),
            .I(N__28845));
    LocalMux I__5019 (
            .O(N__28845),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__5018 (
            .O(N__28842),
            .I(N__28839));
    InMux I__5017 (
            .O(N__28839),
            .I(N__28836));
    LocalMux I__5016 (
            .O(N__28836),
            .I(N__28833));
    Odrv12 I__5015 (
            .O(N__28833),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__5014 (
            .O(N__28830),
            .I(N__28827));
    LocalMux I__5013 (
            .O(N__28827),
            .I(N__28824));
    Odrv4 I__5012 (
            .O(N__28824),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__5011 (
            .O(N__28821),
            .I(N__28818));
    LocalMux I__5010 (
            .O(N__28818),
            .I(N__28815));
    Odrv4 I__5009 (
            .O(N__28815),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__5008 (
            .O(N__28812),
            .I(N__28809));
    InMux I__5007 (
            .O(N__28809),
            .I(N__28806));
    LocalMux I__5006 (
            .O(N__28806),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__5005 (
            .O(N__28803),
            .I(N__28800));
    InMux I__5004 (
            .O(N__28800),
            .I(N__28794));
    InMux I__5003 (
            .O(N__28799),
            .I(N__28794));
    LocalMux I__5002 (
            .O(N__28794),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    InMux I__5001 (
            .O(N__28791),
            .I(N__28788));
    LocalMux I__5000 (
            .O(N__28788),
            .I(N__28785));
    Span4Mux_h I__4999 (
            .O(N__28785),
            .I(N__28782));
    Odrv4 I__4998 (
            .O(N__28782),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__4997 (
            .O(N__28779),
            .I(N__28776));
    InMux I__4996 (
            .O(N__28776),
            .I(N__28773));
    LocalMux I__4995 (
            .O(N__28773),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__4994 (
            .O(N__28770),
            .I(N__28767));
    LocalMux I__4993 (
            .O(N__28767),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__4992 (
            .O(N__28764),
            .I(N__28761));
    InMux I__4991 (
            .O(N__28761),
            .I(N__28758));
    LocalMux I__4990 (
            .O(N__28758),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    InMux I__4989 (
            .O(N__28755),
            .I(N__28752));
    LocalMux I__4988 (
            .O(N__28752),
            .I(N__28749));
    Odrv12 I__4987 (
            .O(N__28749),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__4986 (
            .O(N__28746),
            .I(N__28743));
    InMux I__4985 (
            .O(N__28743),
            .I(N__28740));
    LocalMux I__4984 (
            .O(N__28740),
            .I(N__28737));
    Odrv4 I__4983 (
            .O(N__28737),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__4982 (
            .O(N__28734),
            .I(N__28731));
    LocalMux I__4981 (
            .O(N__28731),
            .I(N__28728));
    Odrv12 I__4980 (
            .O(N__28728),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__4979 (
            .O(N__28725),
            .I(N__28722));
    InMux I__4978 (
            .O(N__28722),
            .I(N__28719));
    LocalMux I__4977 (
            .O(N__28719),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__4976 (
            .O(N__28716),
            .I(N__28713));
    LocalMux I__4975 (
            .O(N__28713),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__4974 (
            .O(N__28710),
            .I(N__28707));
    InMux I__4973 (
            .O(N__28707),
            .I(N__28704));
    LocalMux I__4972 (
            .O(N__28704),
            .I(N__28701));
    Odrv4 I__4971 (
            .O(N__28701),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__4970 (
            .O(N__28698),
            .I(N__28695));
    LocalMux I__4969 (
            .O(N__28695),
            .I(N__28692));
    Span4Mux_h I__4968 (
            .O(N__28692),
            .I(N__28689));
    Odrv4 I__4967 (
            .O(N__28689),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__4966 (
            .O(N__28686),
            .I(N__28683));
    InMux I__4965 (
            .O(N__28683),
            .I(N__28680));
    LocalMux I__4964 (
            .O(N__28680),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__4963 (
            .O(N__28677),
            .I(N__28671));
    InMux I__4962 (
            .O(N__28676),
            .I(N__28664));
    InMux I__4961 (
            .O(N__28675),
            .I(N__28664));
    InMux I__4960 (
            .O(N__28674),
            .I(N__28664));
    LocalMux I__4959 (
            .O(N__28671),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__4958 (
            .O(N__28664),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__4957 (
            .O(N__28659),
            .I(N__28650));
    InMux I__4956 (
            .O(N__28658),
            .I(N__28650));
    InMux I__4955 (
            .O(N__28657),
            .I(N__28650));
    LocalMux I__4954 (
            .O(N__28650),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    CascadeMux I__4953 (
            .O(N__28647),
            .I(N__28642));
    InMux I__4952 (
            .O(N__28646),
            .I(N__28638));
    InMux I__4951 (
            .O(N__28645),
            .I(N__28631));
    InMux I__4950 (
            .O(N__28642),
            .I(N__28631));
    InMux I__4949 (
            .O(N__28641),
            .I(N__28631));
    LocalMux I__4948 (
            .O(N__28638),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    LocalMux I__4947 (
            .O(N__28631),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__4946 (
            .O(N__28626),
            .I(N__28622));
    CascadeMux I__4945 (
            .O(N__28625),
            .I(N__28618));
    InMux I__4944 (
            .O(N__28622),
            .I(N__28611));
    InMux I__4943 (
            .O(N__28621),
            .I(N__28611));
    InMux I__4942 (
            .O(N__28618),
            .I(N__28611));
    LocalMux I__4941 (
            .O(N__28611),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    CascadeMux I__4940 (
            .O(N__28608),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ));
    InMux I__4939 (
            .O(N__28605),
            .I(N__28596));
    InMux I__4938 (
            .O(N__28604),
            .I(N__28596));
    InMux I__4937 (
            .O(N__28603),
            .I(N__28596));
    LocalMux I__4936 (
            .O(N__28596),
            .I(N__28593));
    Odrv4 I__4935 (
            .O(N__28593),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    CascadeMux I__4934 (
            .O(N__28590),
            .I(N__28586));
    InMux I__4933 (
            .O(N__28589),
            .I(N__28578));
    InMux I__4932 (
            .O(N__28586),
            .I(N__28578));
    InMux I__4931 (
            .O(N__28585),
            .I(N__28578));
    LocalMux I__4930 (
            .O(N__28578),
            .I(N__28575));
    Odrv4 I__4929 (
            .O(N__28575),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    CascadeMux I__4928 (
            .O(N__28572),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df30_cascade_ ));
    CascadeMux I__4927 (
            .O(N__28569),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__4926 (
            .O(N__28566),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    CascadeMux I__4925 (
            .O(N__28563),
            .I(N__28559));
    CascadeMux I__4924 (
            .O(N__28562),
            .I(N__28556));
    InMux I__4923 (
            .O(N__28559),
            .I(N__28550));
    InMux I__4922 (
            .O(N__28556),
            .I(N__28550));
    InMux I__4921 (
            .O(N__28555),
            .I(N__28547));
    LocalMux I__4920 (
            .O(N__28550),
            .I(N__28544));
    LocalMux I__4919 (
            .O(N__28547),
            .I(N__28539));
    Span4Mux_v I__4918 (
            .O(N__28544),
            .I(N__28539));
    Odrv4 I__4917 (
            .O(N__28539),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__4916 (
            .O(N__28536),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__4915 (
            .O(N__28533),
            .I(N__28528));
    InMux I__4914 (
            .O(N__28532),
            .I(N__28523));
    InMux I__4913 (
            .O(N__28531),
            .I(N__28523));
    LocalMux I__4912 (
            .O(N__28528),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__4911 (
            .O(N__28523),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__4910 (
            .O(N__28518),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    CascadeMux I__4909 (
            .O(N__28515),
            .I(N__28510));
    InMux I__4908 (
            .O(N__28514),
            .I(N__28507));
    InMux I__4907 (
            .O(N__28513),
            .I(N__28502));
    InMux I__4906 (
            .O(N__28510),
            .I(N__28502));
    LocalMux I__4905 (
            .O(N__28507),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__4904 (
            .O(N__28502),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__4903 (
            .O(N__28497),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__4902 (
            .O(N__28494),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__4901 (
            .O(N__28491),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__4900 (
            .O(N__28488),
            .I(N__28483));
    InMux I__4899 (
            .O(N__28487),
            .I(N__28478));
    InMux I__4898 (
            .O(N__28486),
            .I(N__28478));
    LocalMux I__4897 (
            .O(N__28483),
            .I(N__28474));
    LocalMux I__4896 (
            .O(N__28478),
            .I(N__28471));
    InMux I__4895 (
            .O(N__28477),
            .I(N__28468));
    Span4Mux_v I__4894 (
            .O(N__28474),
            .I(N__28461));
    Span4Mux_v I__4893 (
            .O(N__28471),
            .I(N__28461));
    LocalMux I__4892 (
            .O(N__28468),
            .I(N__28461));
    Span4Mux_h I__4891 (
            .O(N__28461),
            .I(N__28458));
    Span4Mux_v I__4890 (
            .O(N__28458),
            .I(N__28455));
    Odrv4 I__4889 (
            .O(N__28455),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__4888 (
            .O(N__28452),
            .I(N__28449));
    LocalMux I__4887 (
            .O(N__28449),
            .I(N__28446));
    Span4Mux_v I__4886 (
            .O(N__28446),
            .I(N__28441));
    InMux I__4885 (
            .O(N__28445),
            .I(N__28436));
    InMux I__4884 (
            .O(N__28444),
            .I(N__28436));
    Odrv4 I__4883 (
            .O(N__28441),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    LocalMux I__4882 (
            .O(N__28436),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__4881 (
            .O(N__28431),
            .I(N__28424));
    InMux I__4880 (
            .O(N__28430),
            .I(N__28424));
    InMux I__4879 (
            .O(N__28429),
            .I(N__28421));
    LocalMux I__4878 (
            .O(N__28424),
            .I(N__28418));
    LocalMux I__4877 (
            .O(N__28421),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__4876 (
            .O(N__28418),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__4875 (
            .O(N__28413),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    CascadeMux I__4874 (
            .O(N__28410),
            .I(N__28407));
    InMux I__4873 (
            .O(N__28407),
            .I(N__28400));
    InMux I__4872 (
            .O(N__28406),
            .I(N__28400));
    InMux I__4871 (
            .O(N__28405),
            .I(N__28397));
    LocalMux I__4870 (
            .O(N__28400),
            .I(N__28394));
    LocalMux I__4869 (
            .O(N__28397),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv12 I__4868 (
            .O(N__28394),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__4867 (
            .O(N__28389),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    CascadeMux I__4866 (
            .O(N__28386),
            .I(N__28382));
    CascadeMux I__4865 (
            .O(N__28385),
            .I(N__28379));
    InMux I__4864 (
            .O(N__28382),
            .I(N__28376));
    InMux I__4863 (
            .O(N__28379),
            .I(N__28373));
    LocalMux I__4862 (
            .O(N__28376),
            .I(N__28367));
    LocalMux I__4861 (
            .O(N__28373),
            .I(N__28367));
    InMux I__4860 (
            .O(N__28372),
            .I(N__28364));
    Span4Mux_v I__4859 (
            .O(N__28367),
            .I(N__28361));
    LocalMux I__4858 (
            .O(N__28364),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__4857 (
            .O(N__28361),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__4856 (
            .O(N__28356),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__4855 (
            .O(N__28353),
            .I(N__28349));
    InMux I__4854 (
            .O(N__28352),
            .I(N__28345));
    LocalMux I__4853 (
            .O(N__28349),
            .I(N__28342));
    InMux I__4852 (
            .O(N__28348),
            .I(N__28339));
    LocalMux I__4851 (
            .O(N__28345),
            .I(N__28336));
    Span4Mux_h I__4850 (
            .O(N__28342),
            .I(N__28333));
    LocalMux I__4849 (
            .O(N__28339),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__4848 (
            .O(N__28336),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__4847 (
            .O(N__28333),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__4846 (
            .O(N__28326),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__4845 (
            .O(N__28323),
            .I(N__28319));
    InMux I__4844 (
            .O(N__28322),
            .I(N__28313));
    InMux I__4843 (
            .O(N__28319),
            .I(N__28313));
    InMux I__4842 (
            .O(N__28318),
            .I(N__28310));
    LocalMux I__4841 (
            .O(N__28313),
            .I(N__28307));
    LocalMux I__4840 (
            .O(N__28310),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__4839 (
            .O(N__28307),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__4838 (
            .O(N__28302),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    CascadeMux I__4837 (
            .O(N__28299),
            .I(N__28296));
    InMux I__4836 (
            .O(N__28296),
            .I(N__28291));
    InMux I__4835 (
            .O(N__28295),
            .I(N__28288));
    InMux I__4834 (
            .O(N__28294),
            .I(N__28285));
    LocalMux I__4833 (
            .O(N__28291),
            .I(N__28280));
    LocalMux I__4832 (
            .O(N__28288),
            .I(N__28280));
    LocalMux I__4831 (
            .O(N__28285),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__4830 (
            .O(N__28280),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__4829 (
            .O(N__28275),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__4828 (
            .O(N__28272),
            .I(N__28265));
    InMux I__4827 (
            .O(N__28271),
            .I(N__28265));
    InMux I__4826 (
            .O(N__28270),
            .I(N__28262));
    LocalMux I__4825 (
            .O(N__28265),
            .I(N__28259));
    LocalMux I__4824 (
            .O(N__28262),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__4823 (
            .O(N__28259),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__4822 (
            .O(N__28254),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    CascadeMux I__4821 (
            .O(N__28251),
            .I(N__28247));
    InMux I__4820 (
            .O(N__28250),
            .I(N__28241));
    InMux I__4819 (
            .O(N__28247),
            .I(N__28241));
    InMux I__4818 (
            .O(N__28246),
            .I(N__28238));
    LocalMux I__4817 (
            .O(N__28241),
            .I(N__28235));
    LocalMux I__4816 (
            .O(N__28238),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__4815 (
            .O(N__28235),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__4814 (
            .O(N__28230),
            .I(bfn_11_8_0_));
    InMux I__4813 (
            .O(N__28227),
            .I(N__28220));
    InMux I__4812 (
            .O(N__28226),
            .I(N__28220));
    InMux I__4811 (
            .O(N__28225),
            .I(N__28217));
    LocalMux I__4810 (
            .O(N__28220),
            .I(N__28214));
    LocalMux I__4809 (
            .O(N__28217),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    Odrv4 I__4808 (
            .O(N__28214),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__4807 (
            .O(N__28209),
            .I(bfn_11_6_0_));
    InMux I__4806 (
            .O(N__28206),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__4805 (
            .O(N__28203),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__4804 (
            .O(N__28200),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__4803 (
            .O(N__28197),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__4802 (
            .O(N__28194),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__4801 (
            .O(N__28191),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__4800 (
            .O(N__28188),
            .I(N__28181));
    InMux I__4799 (
            .O(N__28187),
            .I(N__28181));
    InMux I__4798 (
            .O(N__28186),
            .I(N__28178));
    LocalMux I__4797 (
            .O(N__28181),
            .I(N__28175));
    LocalMux I__4796 (
            .O(N__28178),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__4795 (
            .O(N__28175),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__4794 (
            .O(N__28170),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    CascadeMux I__4793 (
            .O(N__28167),
            .I(N__28162));
    InMux I__4792 (
            .O(N__28166),
            .I(N__28159));
    InMux I__4791 (
            .O(N__28165),
            .I(N__28154));
    InMux I__4790 (
            .O(N__28162),
            .I(N__28154));
    LocalMux I__4789 (
            .O(N__28159),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__4788 (
            .O(N__28154),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__4787 (
            .O(N__28149),
            .I(bfn_11_7_0_));
    CascadeMux I__4786 (
            .O(N__28146),
            .I(N__28143));
    InMux I__4785 (
            .O(N__28143),
            .I(N__28136));
    InMux I__4784 (
            .O(N__28142),
            .I(N__28136));
    InMux I__4783 (
            .O(N__28141),
            .I(N__28133));
    LocalMux I__4782 (
            .O(N__28136),
            .I(N__28130));
    LocalMux I__4781 (
            .O(N__28133),
            .I(N__28125));
    Span4Mux_h I__4780 (
            .O(N__28130),
            .I(N__28125));
    Span4Mux_v I__4779 (
            .O(N__28125),
            .I(N__28122));
    Span4Mux_v I__4778 (
            .O(N__28122),
            .I(N__28119));
    Odrv4 I__4777 (
            .O(N__28119),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__4776 (
            .O(N__28116),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__4775 (
            .O(N__28113),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__4774 (
            .O(N__28110),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__4773 (
            .O(N__28107),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__4772 (
            .O(N__28104),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__4771 (
            .O(N__28101),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__4770 (
            .O(N__28098),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    CascadeMux I__4769 (
            .O(N__28095),
            .I(N__28092));
    InMux I__4768 (
            .O(N__28092),
            .I(N__28089));
    LocalMux I__4767 (
            .O(N__28089),
            .I(N__28086));
    Span4Mux_v I__4766 (
            .O(N__28086),
            .I(N__28083));
    Span4Mux_h I__4765 (
            .O(N__28083),
            .I(N__28080));
    Span4Mux_h I__4764 (
            .O(N__28080),
            .I(N__28077));
    Span4Mux_h I__4763 (
            .O(N__28077),
            .I(N__28074));
    Odrv4 I__4762 (
            .O(N__28074),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    InMux I__4761 (
            .O(N__28071),
            .I(N__28068));
    LocalMux I__4760 (
            .O(N__28068),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ));
    InMux I__4759 (
            .O(N__28065),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    CascadeMux I__4758 (
            .O(N__28062),
            .I(N__28059));
    InMux I__4757 (
            .O(N__28059),
            .I(N__28056));
    LocalMux I__4756 (
            .O(N__28056),
            .I(N__28053));
    Span4Mux_v I__4755 (
            .O(N__28053),
            .I(N__28050));
    Sp12to4 I__4754 (
            .O(N__28050),
            .I(N__28047));
    Span12Mux_h I__4753 (
            .O(N__28047),
            .I(N__28044));
    Odrv12 I__4752 (
            .O(N__28044),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__4751 (
            .O(N__28041),
            .I(N__28038));
    LocalMux I__4750 (
            .O(N__28038),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ));
    InMux I__4749 (
            .O(N__28035),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    CascadeMux I__4748 (
            .O(N__28032),
            .I(N__28029));
    InMux I__4747 (
            .O(N__28029),
            .I(N__28026));
    LocalMux I__4746 (
            .O(N__28026),
            .I(N__28023));
    Span12Mux_h I__4745 (
            .O(N__28023),
            .I(N__28020));
    Span12Mux_h I__4744 (
            .O(N__28020),
            .I(N__28017));
    Odrv12 I__4743 (
            .O(N__28017),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__4742 (
            .O(N__28014),
            .I(N__28011));
    LocalMux I__4741 (
            .O(N__28011),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ));
    InMux I__4740 (
            .O(N__28008),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    CascadeMux I__4739 (
            .O(N__28005),
            .I(N__28002));
    InMux I__4738 (
            .O(N__28002),
            .I(N__27999));
    LocalMux I__4737 (
            .O(N__27999),
            .I(N__27996));
    Span4Mux_v I__4736 (
            .O(N__27996),
            .I(N__27993));
    Sp12to4 I__4735 (
            .O(N__27993),
            .I(N__27990));
    Span12Mux_h I__4734 (
            .O(N__27990),
            .I(N__27987));
    Odrv12 I__4733 (
            .O(N__27987),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__4732 (
            .O(N__27984),
            .I(N__27981));
    LocalMux I__4731 (
            .O(N__27981),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ));
    InMux I__4730 (
            .O(N__27978),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    CascadeMux I__4729 (
            .O(N__27975),
            .I(N__27972));
    InMux I__4728 (
            .O(N__27972),
            .I(N__27969));
    LocalMux I__4727 (
            .O(N__27969),
            .I(N__27966));
    Span4Mux_v I__4726 (
            .O(N__27966),
            .I(N__27963));
    Sp12to4 I__4725 (
            .O(N__27963),
            .I(N__27960));
    Span12Mux_h I__4724 (
            .O(N__27960),
            .I(N__27957));
    Odrv12 I__4723 (
            .O(N__27957),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    InMux I__4722 (
            .O(N__27954),
            .I(N__27951));
    LocalMux I__4721 (
            .O(N__27951),
            .I(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ));
    InMux I__4720 (
            .O(N__27948),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    CascadeMux I__4719 (
            .O(N__27945),
            .I(N__27942));
    InMux I__4718 (
            .O(N__27942),
            .I(N__27939));
    LocalMux I__4717 (
            .O(N__27939),
            .I(N__27936));
    Span4Mux_v I__4716 (
            .O(N__27936),
            .I(N__27933));
    Span4Mux_h I__4715 (
            .O(N__27933),
            .I(N__27930));
    Sp12to4 I__4714 (
            .O(N__27930),
            .I(N__27927));
    Odrv12 I__4713 (
            .O(N__27927),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__4712 (
            .O(N__27924),
            .I(N__27921));
    LocalMux I__4711 (
            .O(N__27921),
            .I(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ));
    InMux I__4710 (
            .O(N__27918),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    InMux I__4709 (
            .O(N__27915),
            .I(N__27903));
    InMux I__4708 (
            .O(N__27914),
            .I(N__27903));
    InMux I__4707 (
            .O(N__27913),
            .I(N__27896));
    InMux I__4706 (
            .O(N__27912),
            .I(N__27896));
    InMux I__4705 (
            .O(N__27911),
            .I(N__27896));
    InMux I__4704 (
            .O(N__27910),
            .I(N__27889));
    InMux I__4703 (
            .O(N__27909),
            .I(N__27889));
    InMux I__4702 (
            .O(N__27908),
            .I(N__27889));
    LocalMux I__4701 (
            .O(N__27903),
            .I(N__27886));
    LocalMux I__4700 (
            .O(N__27896),
            .I(N__27881));
    LocalMux I__4699 (
            .O(N__27889),
            .I(N__27881));
    Span12Mux_h I__4698 (
            .O(N__27886),
            .I(N__27878));
    Span12Mux_h I__4697 (
            .O(N__27881),
            .I(N__27875));
    Odrv12 I__4696 (
            .O(N__27878),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    Odrv12 I__4695 (
            .O(N__27875),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    CascadeMux I__4694 (
            .O(N__27870),
            .I(N__27867));
    InMux I__4693 (
            .O(N__27867),
            .I(N__27864));
    LocalMux I__4692 (
            .O(N__27864),
            .I(N__27861));
    Odrv12 I__4691 (
            .O(N__27861),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    InMux I__4690 (
            .O(N__27858),
            .I(N__27855));
    LocalMux I__4689 (
            .O(N__27855),
            .I(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ));
    InMux I__4688 (
            .O(N__27852),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__4687 (
            .O(N__27849),
            .I(N__27846));
    LocalMux I__4686 (
            .O(N__27846),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__4685 (
            .O(N__27843),
            .I(N__27840));
    LocalMux I__4684 (
            .O(N__27840),
            .I(N__27837));
    Odrv12 I__4683 (
            .O(N__27837),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__4682 (
            .O(N__27834),
            .I(bfn_10_28_0_));
    InMux I__4681 (
            .O(N__27831),
            .I(N__27828));
    LocalMux I__4680 (
            .O(N__27828),
            .I(N__27825));
    Span4Mux_v I__4679 (
            .O(N__27825),
            .I(N__27822));
    Sp12to4 I__4678 (
            .O(N__27822),
            .I(N__27819));
    Span12Mux_h I__4677 (
            .O(N__27819),
            .I(N__27816));
    Odrv12 I__4676 (
            .O(N__27816),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__4675 (
            .O(N__27813),
            .I(N__27810));
    InMux I__4674 (
            .O(N__27810),
            .I(N__27807));
    LocalMux I__4673 (
            .O(N__27807),
            .I(N__27804));
    Span12Mux_h I__4672 (
            .O(N__27804),
            .I(N__27801));
    Odrv12 I__4671 (
            .O(N__27801),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__4670 (
            .O(N__27798),
            .I(N__27795));
    LocalMux I__4669 (
            .O(N__27795),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ));
    InMux I__4668 (
            .O(N__27792),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__4667 (
            .O(N__27789),
            .I(N__27786));
    LocalMux I__4666 (
            .O(N__27786),
            .I(N__27783));
    Span12Mux_h I__4665 (
            .O(N__27783),
            .I(N__27780));
    Span12Mux_h I__4664 (
            .O(N__27780),
            .I(N__27777));
    Odrv12 I__4663 (
            .O(N__27777),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__4662 (
            .O(N__27774),
            .I(N__27771));
    InMux I__4661 (
            .O(N__27771),
            .I(N__27768));
    LocalMux I__4660 (
            .O(N__27768),
            .I(N__27765));
    Span4Mux_h I__4659 (
            .O(N__27765),
            .I(N__27762));
    Span4Mux_h I__4658 (
            .O(N__27762),
            .I(N__27759));
    Span4Mux_h I__4657 (
            .O(N__27759),
            .I(N__27756));
    Odrv4 I__4656 (
            .O(N__27756),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    CascadeMux I__4655 (
            .O(N__27753),
            .I(N__27750));
    InMux I__4654 (
            .O(N__27750),
            .I(N__27747));
    LocalMux I__4653 (
            .O(N__27747),
            .I(N__27744));
    Odrv4 I__4652 (
            .O(N__27744),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ));
    InMux I__4651 (
            .O(N__27741),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__4650 (
            .O(N__27738),
            .I(N__27735));
    LocalMux I__4649 (
            .O(N__27735),
            .I(N__27732));
    Span4Mux_v I__4648 (
            .O(N__27732),
            .I(N__27729));
    Sp12to4 I__4647 (
            .O(N__27729),
            .I(N__27726));
    Span12Mux_h I__4646 (
            .O(N__27726),
            .I(N__27723));
    Odrv12 I__4645 (
            .O(N__27723),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    CascadeMux I__4644 (
            .O(N__27720),
            .I(N__27717));
    InMux I__4643 (
            .O(N__27717),
            .I(N__27714));
    LocalMux I__4642 (
            .O(N__27714),
            .I(N__27711));
    Span4Mux_h I__4641 (
            .O(N__27711),
            .I(N__27708));
    Span4Mux_h I__4640 (
            .O(N__27708),
            .I(N__27705));
    Span4Mux_h I__4639 (
            .O(N__27705),
            .I(N__27702));
    Odrv4 I__4638 (
            .O(N__27702),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__4637 (
            .O(N__27699),
            .I(N__27696));
    LocalMux I__4636 (
            .O(N__27696),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ));
    InMux I__4635 (
            .O(N__27693),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__4634 (
            .O(N__27690),
            .I(N__27687));
    LocalMux I__4633 (
            .O(N__27687),
            .I(N__27684));
    Span4Mux_v I__4632 (
            .O(N__27684),
            .I(N__27681));
    Sp12to4 I__4631 (
            .O(N__27681),
            .I(N__27678));
    Span12Mux_h I__4630 (
            .O(N__27678),
            .I(N__27675));
    Odrv12 I__4629 (
            .O(N__27675),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__4628 (
            .O(N__27672),
            .I(N__27669));
    InMux I__4627 (
            .O(N__27669),
            .I(N__27666));
    LocalMux I__4626 (
            .O(N__27666),
            .I(N__27663));
    Span4Mux_v I__4625 (
            .O(N__27663),
            .I(N__27660));
    Span4Mux_h I__4624 (
            .O(N__27660),
            .I(N__27657));
    Span4Mux_h I__4623 (
            .O(N__27657),
            .I(N__27654));
    Odrv4 I__4622 (
            .O(N__27654),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    InMux I__4621 (
            .O(N__27651),
            .I(N__27648));
    LocalMux I__4620 (
            .O(N__27648),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ));
    InMux I__4619 (
            .O(N__27645),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__4618 (
            .O(N__27642),
            .I(N__27639));
    LocalMux I__4617 (
            .O(N__27639),
            .I(N__27636));
    Span4Mux_v I__4616 (
            .O(N__27636),
            .I(N__27633));
    Span4Mux_h I__4615 (
            .O(N__27633),
            .I(N__27630));
    Sp12to4 I__4614 (
            .O(N__27630),
            .I(N__27627));
    Odrv12 I__4613 (
            .O(N__27627),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    CascadeMux I__4612 (
            .O(N__27624),
            .I(N__27621));
    InMux I__4611 (
            .O(N__27621),
            .I(N__27618));
    LocalMux I__4610 (
            .O(N__27618),
            .I(N__27615));
    Sp12to4 I__4609 (
            .O(N__27615),
            .I(N__27612));
    Span12Mux_s5_v I__4608 (
            .O(N__27612),
            .I(N__27609));
    Odrv12 I__4607 (
            .O(N__27609),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    InMux I__4606 (
            .O(N__27606),
            .I(N__27603));
    LocalMux I__4605 (
            .O(N__27603),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ));
    InMux I__4604 (
            .O(N__27600),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__4603 (
            .O(N__27597),
            .I(N__27594));
    LocalMux I__4602 (
            .O(N__27594),
            .I(N__27591));
    Span12Mux_s5_v I__4601 (
            .O(N__27591),
            .I(N__27588));
    Odrv12 I__4600 (
            .O(N__27588),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    CascadeMux I__4599 (
            .O(N__27585),
            .I(N__27582));
    InMux I__4598 (
            .O(N__27582),
            .I(N__27579));
    LocalMux I__4597 (
            .O(N__27579),
            .I(N__27576));
    Span12Mux_s7_v I__4596 (
            .O(N__27576),
            .I(N__27573));
    Span12Mux_h I__4595 (
            .O(N__27573),
            .I(N__27570));
    Odrv12 I__4594 (
            .O(N__27570),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    InMux I__4593 (
            .O(N__27567),
            .I(N__27564));
    LocalMux I__4592 (
            .O(N__27564),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ));
    InMux I__4591 (
            .O(N__27561),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__4590 (
            .O(N__27558),
            .I(N__27555));
    LocalMux I__4589 (
            .O(N__27555),
            .I(N__27552));
    Span4Mux_v I__4588 (
            .O(N__27552),
            .I(N__27549));
    Sp12to4 I__4587 (
            .O(N__27549),
            .I(N__27546));
    Odrv12 I__4586 (
            .O(N__27546),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    CascadeMux I__4585 (
            .O(N__27543),
            .I(N__27540));
    InMux I__4584 (
            .O(N__27540),
            .I(N__27537));
    LocalMux I__4583 (
            .O(N__27537),
            .I(N__27534));
    Span4Mux_v I__4582 (
            .O(N__27534),
            .I(N__27531));
    Sp12to4 I__4581 (
            .O(N__27531),
            .I(N__27528));
    Span12Mux_h I__4580 (
            .O(N__27528),
            .I(N__27525));
    Odrv12 I__4579 (
            .O(N__27525),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    InMux I__4578 (
            .O(N__27522),
            .I(N__27519));
    LocalMux I__4577 (
            .O(N__27519),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ));
    InMux I__4576 (
            .O(N__27516),
            .I(bfn_10_27_0_));
    InMux I__4575 (
            .O(N__27513),
            .I(N__27510));
    LocalMux I__4574 (
            .O(N__27510),
            .I(N__27507));
    Span4Mux_h I__4573 (
            .O(N__27507),
            .I(N__27504));
    Span4Mux_h I__4572 (
            .O(N__27504),
            .I(N__27501));
    Span4Mux_h I__4571 (
            .O(N__27501),
            .I(N__27498));
    Odrv4 I__4570 (
            .O(N__27498),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    InMux I__4569 (
            .O(N__27495),
            .I(N__27489));
    InMux I__4568 (
            .O(N__27494),
            .I(N__27489));
    LocalMux I__4567 (
            .O(N__27489),
            .I(N__27486));
    Span12Mux_v I__4566 (
            .O(N__27486),
            .I(N__27483));
    Span12Mux_h I__4565 (
            .O(N__27483),
            .I(N__27480));
    Odrv12 I__4564 (
            .O(N__27480),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    InMux I__4563 (
            .O(N__27477),
            .I(N__27474));
    LocalMux I__4562 (
            .O(N__27474),
            .I(N__27471));
    Span4Mux_v I__4561 (
            .O(N__27471),
            .I(N__27468));
    Sp12to4 I__4560 (
            .O(N__27468),
            .I(N__27465));
    Span12Mux_h I__4559 (
            .O(N__27465),
            .I(N__27462));
    Odrv12 I__4558 (
            .O(N__27462),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__4557 (
            .O(N__27459),
            .I(N__27456));
    LocalMux I__4556 (
            .O(N__27456),
            .I(N__27453));
    Span4Mux_h I__4555 (
            .O(N__27453),
            .I(N__27450));
    Odrv4 I__4554 (
            .O(N__27450),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__4553 (
            .O(N__27447),
            .I(N__27443));
    InMux I__4552 (
            .O(N__27446),
            .I(N__27440));
    LocalMux I__4551 (
            .O(N__27443),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    LocalMux I__4550 (
            .O(N__27440),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    InMux I__4549 (
            .O(N__27435),
            .I(N__27432));
    LocalMux I__4548 (
            .O(N__27432),
            .I(N__27428));
    InMux I__4547 (
            .O(N__27431),
            .I(N__27424));
    Span4Mux_h I__4546 (
            .O(N__27428),
            .I(N__27421));
    InMux I__4545 (
            .O(N__27427),
            .I(N__27418));
    LocalMux I__4544 (
            .O(N__27424),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    Odrv4 I__4543 (
            .O(N__27421),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    LocalMux I__4542 (
            .O(N__27418),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__4541 (
            .O(N__27411),
            .I(N__27408));
    LocalMux I__4540 (
            .O(N__27408),
            .I(N__27405));
    Span4Mux_h I__4539 (
            .O(N__27405),
            .I(N__27402));
    Odrv4 I__4538 (
            .O(N__27402),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    CascadeMux I__4537 (
            .O(N__27399),
            .I(N__27396));
    InMux I__4536 (
            .O(N__27396),
            .I(N__27393));
    LocalMux I__4535 (
            .O(N__27393),
            .I(N__27389));
    InMux I__4534 (
            .O(N__27392),
            .I(N__27385));
    Span4Mux_v I__4533 (
            .O(N__27389),
            .I(N__27382));
    InMux I__4532 (
            .O(N__27388),
            .I(N__27379));
    LocalMux I__4531 (
            .O(N__27385),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    Odrv4 I__4530 (
            .O(N__27382),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__4529 (
            .O(N__27379),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    InMux I__4528 (
            .O(N__27372),
            .I(N__27368));
    InMux I__4527 (
            .O(N__27371),
            .I(N__27365));
    LocalMux I__4526 (
            .O(N__27368),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    LocalMux I__4525 (
            .O(N__27365),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    InMux I__4524 (
            .O(N__27360),
            .I(N__27357));
    LocalMux I__4523 (
            .O(N__27357),
            .I(N__27354));
    Span4Mux_h I__4522 (
            .O(N__27354),
            .I(N__27351));
    Odrv4 I__4521 (
            .O(N__27351),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    CascadeMux I__4520 (
            .O(N__27348),
            .I(N__27345));
    InMux I__4519 (
            .O(N__27345),
            .I(N__27341));
    InMux I__4518 (
            .O(N__27344),
            .I(N__27338));
    LocalMux I__4517 (
            .O(N__27341),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    LocalMux I__4516 (
            .O(N__27338),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    InMux I__4515 (
            .O(N__27333),
            .I(N__27330));
    LocalMux I__4514 (
            .O(N__27330),
            .I(N__27326));
    InMux I__4513 (
            .O(N__27329),
            .I(N__27322));
    Span4Mux_h I__4512 (
            .O(N__27326),
            .I(N__27319));
    InMux I__4511 (
            .O(N__27325),
            .I(N__27316));
    LocalMux I__4510 (
            .O(N__27322),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__4509 (
            .O(N__27319),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    LocalMux I__4508 (
            .O(N__27316),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__4507 (
            .O(N__27309),
            .I(N__27304));
    InMux I__4506 (
            .O(N__27308),
            .I(N__27301));
    InMux I__4505 (
            .O(N__27307),
            .I(N__27298));
    LocalMux I__4504 (
            .O(N__27304),
            .I(N__27295));
    LocalMux I__4503 (
            .O(N__27301),
            .I(N__27292));
    LocalMux I__4502 (
            .O(N__27298),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv12 I__4501 (
            .O(N__27295),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__4500 (
            .O(N__27292),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    InMux I__4499 (
            .O(N__27285),
            .I(N__27282));
    LocalMux I__4498 (
            .O(N__27282),
            .I(N__27279));
    Span4Mux_v I__4497 (
            .O(N__27279),
            .I(N__27276));
    Odrv4 I__4496 (
            .O(N__27276),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    InMux I__4495 (
            .O(N__27273),
            .I(N__27270));
    LocalMux I__4494 (
            .O(N__27270),
            .I(N__27266));
    InMux I__4493 (
            .O(N__27269),
            .I(N__27263));
    Span4Mux_h I__4492 (
            .O(N__27266),
            .I(N__27258));
    LocalMux I__4491 (
            .O(N__27263),
            .I(N__27258));
    Span4Mux_h I__4490 (
            .O(N__27258),
            .I(N__27255));
    Span4Mux_h I__4489 (
            .O(N__27255),
            .I(N__27252));
    Odrv4 I__4488 (
            .O(N__27252),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__4487 (
            .O(N__27249),
            .I(N__27245));
    InMux I__4486 (
            .O(N__27248),
            .I(N__27242));
    LocalMux I__4485 (
            .O(N__27245),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    LocalMux I__4484 (
            .O(N__27242),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    CascadeMux I__4483 (
            .O(N__27237),
            .I(N__27234));
    InMux I__4482 (
            .O(N__27234),
            .I(N__27231));
    LocalMux I__4481 (
            .O(N__27231),
            .I(N__27227));
    InMux I__4480 (
            .O(N__27230),
            .I(N__27223));
    Span4Mux_h I__4479 (
            .O(N__27227),
            .I(N__27220));
    InMux I__4478 (
            .O(N__27226),
            .I(N__27217));
    LocalMux I__4477 (
            .O(N__27223),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    Odrv4 I__4476 (
            .O(N__27220),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    LocalMux I__4475 (
            .O(N__27217),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    InMux I__4474 (
            .O(N__27210),
            .I(N__27207));
    LocalMux I__4473 (
            .O(N__27207),
            .I(N__27204));
    Span4Mux_h I__4472 (
            .O(N__27204),
            .I(N__27201));
    Odrv4 I__4471 (
            .O(N__27201),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    InMux I__4470 (
            .O(N__27198),
            .I(N__27195));
    LocalMux I__4469 (
            .O(N__27195),
            .I(N__27192));
    Span4Mux_v I__4468 (
            .O(N__27192),
            .I(N__27189));
    Sp12to4 I__4467 (
            .O(N__27189),
            .I(N__27186));
    Span12Mux_h I__4466 (
            .O(N__27186),
            .I(N__27183));
    Odrv12 I__4465 (
            .O(N__27183),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__4464 (
            .O(N__27180),
            .I(N__27177));
    InMux I__4463 (
            .O(N__27177),
            .I(N__27174));
    LocalMux I__4462 (
            .O(N__27174),
            .I(N__27171));
    Span4Mux_h I__4461 (
            .O(N__27171),
            .I(N__27168));
    Span4Mux_h I__4460 (
            .O(N__27168),
            .I(N__27165));
    Span4Mux_h I__4459 (
            .O(N__27165),
            .I(N__27162));
    Odrv4 I__4458 (
            .O(N__27162),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__4457 (
            .O(N__27159),
            .I(N__27156));
    LocalMux I__4456 (
            .O(N__27156),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__4455 (
            .O(N__27153),
            .I(N__27150));
    LocalMux I__4454 (
            .O(N__27150),
            .I(N__27147));
    Span4Mux_v I__4453 (
            .O(N__27147),
            .I(N__27144));
    Sp12to4 I__4452 (
            .O(N__27144),
            .I(N__27141));
    Span12Mux_h I__4451 (
            .O(N__27141),
            .I(N__27138));
    Odrv12 I__4450 (
            .O(N__27138),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__4449 (
            .O(N__27135),
            .I(N__27132));
    InMux I__4448 (
            .O(N__27132),
            .I(N__27129));
    LocalMux I__4447 (
            .O(N__27129),
            .I(N__27126));
    Span4Mux_h I__4446 (
            .O(N__27126),
            .I(N__27123));
    Span4Mux_h I__4445 (
            .O(N__27123),
            .I(N__27120));
    Span4Mux_h I__4444 (
            .O(N__27120),
            .I(N__27117));
    Odrv4 I__4443 (
            .O(N__27117),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    CascadeMux I__4442 (
            .O(N__27114),
            .I(N__27111));
    InMux I__4441 (
            .O(N__27111),
            .I(N__27108));
    LocalMux I__4440 (
            .O(N__27108),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ));
    InMux I__4439 (
            .O(N__27105),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__4438 (
            .O(N__27102),
            .I(N__27098));
    InMux I__4437 (
            .O(N__27101),
            .I(N__27094));
    LocalMux I__4436 (
            .O(N__27098),
            .I(N__27091));
    InMux I__4435 (
            .O(N__27097),
            .I(N__27088));
    LocalMux I__4434 (
            .O(N__27094),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv12 I__4433 (
            .O(N__27091),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    LocalMux I__4432 (
            .O(N__27088),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    InMux I__4431 (
            .O(N__27081),
            .I(N__27075));
    CascadeMux I__4430 (
            .O(N__27080),
            .I(N__27072));
    InMux I__4429 (
            .O(N__27079),
            .I(N__27069));
    InMux I__4428 (
            .O(N__27078),
            .I(N__27066));
    LocalMux I__4427 (
            .O(N__27075),
            .I(N__27063));
    InMux I__4426 (
            .O(N__27072),
            .I(N__27060));
    LocalMux I__4425 (
            .O(N__27069),
            .I(N__27057));
    LocalMux I__4424 (
            .O(N__27066),
            .I(N__27054));
    Span4Mux_h I__4423 (
            .O(N__27063),
            .I(N__27051));
    LocalMux I__4422 (
            .O(N__27060),
            .I(N__27048));
    Span12Mux_s11_v I__4421 (
            .O(N__27057),
            .I(N__27045));
    Span4Mux_h I__4420 (
            .O(N__27054),
            .I(N__27038));
    Span4Mux_v I__4419 (
            .O(N__27051),
            .I(N__27038));
    Span4Mux_h I__4418 (
            .O(N__27048),
            .I(N__27038));
    Odrv12 I__4417 (
            .O(N__27045),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__4416 (
            .O(N__27038),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    CascadeMux I__4415 (
            .O(N__27033),
            .I(N__27030));
    InMux I__4414 (
            .O(N__27030),
            .I(N__27024));
    InMux I__4413 (
            .O(N__27029),
            .I(N__27024));
    LocalMux I__4412 (
            .O(N__27024),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ));
    CEMux I__4411 (
            .O(N__27021),
            .I(N__27000));
    CEMux I__4410 (
            .O(N__27020),
            .I(N__27000));
    CEMux I__4409 (
            .O(N__27019),
            .I(N__27000));
    CEMux I__4408 (
            .O(N__27018),
            .I(N__27000));
    CEMux I__4407 (
            .O(N__27017),
            .I(N__27000));
    CEMux I__4406 (
            .O(N__27016),
            .I(N__27000));
    CEMux I__4405 (
            .O(N__27015),
            .I(N__27000));
    GlobalMux I__4404 (
            .O(N__27000),
            .I(N__26997));
    gio2CtrlBuf I__4403 (
            .O(N__26997),
            .I(\phase_controller_inst2.stoper_hc.un1_start_g ));
    InMux I__4402 (
            .O(N__26994),
            .I(N__26990));
    InMux I__4401 (
            .O(N__26993),
            .I(N__26987));
    LocalMux I__4400 (
            .O(N__26990),
            .I(N__26984));
    LocalMux I__4399 (
            .O(N__26987),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    Odrv4 I__4398 (
            .O(N__26984),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    InMux I__4397 (
            .O(N__26979),
            .I(N__26975));
    InMux I__4396 (
            .O(N__26978),
            .I(N__26972));
    LocalMux I__4395 (
            .O(N__26975),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    LocalMux I__4394 (
            .O(N__26972),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    InMux I__4393 (
            .O(N__26967),
            .I(N__26961));
    InMux I__4392 (
            .O(N__26966),
            .I(N__26954));
    InMux I__4391 (
            .O(N__26965),
            .I(N__26954));
    InMux I__4390 (
            .O(N__26964),
            .I(N__26954));
    LocalMux I__4389 (
            .O(N__26961),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__4388 (
            .O(N__26954),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__4387 (
            .O(N__26949),
            .I(N__26946));
    LocalMux I__4386 (
            .O(N__26946),
            .I(N__26943));
    Span4Mux_h I__4385 (
            .O(N__26943),
            .I(N__26940));
    Odrv4 I__4384 (
            .O(N__26940),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__4383 (
            .O(N__26937),
            .I(N__26934));
    LocalMux I__4382 (
            .O(N__26934),
            .I(N__26931));
    Span4Mux_h I__4381 (
            .O(N__26931),
            .I(N__26928));
    Odrv4 I__4380 (
            .O(N__26928),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__4379 (
            .O(N__26925),
            .I(N__26922));
    LocalMux I__4378 (
            .O(N__26922),
            .I(N__26919));
    Span4Mux_h I__4377 (
            .O(N__26919),
            .I(N__26916));
    Odrv4 I__4376 (
            .O(N__26916),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__4375 (
            .O(N__26913),
            .I(N__26905));
    InMux I__4374 (
            .O(N__26912),
            .I(N__26893));
    InMux I__4373 (
            .O(N__26911),
            .I(N__26893));
    InMux I__4372 (
            .O(N__26910),
            .I(N__26893));
    InMux I__4371 (
            .O(N__26909),
            .I(N__26893));
    InMux I__4370 (
            .O(N__26908),
            .I(N__26890));
    LocalMux I__4369 (
            .O(N__26905),
            .I(N__26887));
    CascadeMux I__4368 (
            .O(N__26904),
            .I(N__26883));
    InMux I__4367 (
            .O(N__26903),
            .I(N__26878));
    InMux I__4366 (
            .O(N__26902),
            .I(N__26878));
    LocalMux I__4365 (
            .O(N__26893),
            .I(N__26873));
    LocalMux I__4364 (
            .O(N__26890),
            .I(N__26873));
    Span4Mux_h I__4363 (
            .O(N__26887),
            .I(N__26870));
    InMux I__4362 (
            .O(N__26886),
            .I(N__26865));
    InMux I__4361 (
            .O(N__26883),
            .I(N__26865));
    LocalMux I__4360 (
            .O(N__26878),
            .I(N__26862));
    Span4Mux_v I__4359 (
            .O(N__26873),
            .I(N__26859));
    Span4Mux_h I__4358 (
            .O(N__26870),
            .I(N__26854));
    LocalMux I__4357 (
            .O(N__26865),
            .I(N__26854));
    Span4Mux_h I__4356 (
            .O(N__26862),
            .I(N__26851));
    Odrv4 I__4355 (
            .O(N__26859),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__4354 (
            .O(N__26854),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__4353 (
            .O(N__26851),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__4352 (
            .O(N__26844),
            .I(N__26838));
    InMux I__4351 (
            .O(N__26843),
            .I(N__26838));
    LocalMux I__4350 (
            .O(N__26838),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ));
    InMux I__4349 (
            .O(N__26835),
            .I(N__26832));
    LocalMux I__4348 (
            .O(N__26832),
            .I(N__26828));
    InMux I__4347 (
            .O(N__26831),
            .I(N__26824));
    Span4Mux_h I__4346 (
            .O(N__26828),
            .I(N__26821));
    InMux I__4345 (
            .O(N__26827),
            .I(N__26818));
    LocalMux I__4344 (
            .O(N__26824),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    Odrv4 I__4343 (
            .O(N__26821),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    LocalMux I__4342 (
            .O(N__26818),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    InMux I__4341 (
            .O(N__26811),
            .I(N__26808));
    LocalMux I__4340 (
            .O(N__26808),
            .I(N__26802));
    InMux I__4339 (
            .O(N__26807),
            .I(N__26799));
    InMux I__4338 (
            .O(N__26806),
            .I(N__26794));
    InMux I__4337 (
            .O(N__26805),
            .I(N__26794));
    Span4Mux_v I__4336 (
            .O(N__26802),
            .I(N__26789));
    LocalMux I__4335 (
            .O(N__26799),
            .I(N__26789));
    LocalMux I__4334 (
            .O(N__26794),
            .I(N__26786));
    Span4Mux_v I__4333 (
            .O(N__26789),
            .I(N__26783));
    Span4Mux_h I__4332 (
            .O(N__26786),
            .I(N__26780));
    Odrv4 I__4331 (
            .O(N__26783),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    Odrv4 I__4330 (
            .O(N__26780),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    CascadeMux I__4329 (
            .O(N__26775),
            .I(N__26772));
    InMux I__4328 (
            .O(N__26772),
            .I(N__26766));
    InMux I__4327 (
            .O(N__26771),
            .I(N__26766));
    LocalMux I__4326 (
            .O(N__26766),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ));
    InMux I__4325 (
            .O(N__26763),
            .I(N__26759));
    InMux I__4324 (
            .O(N__26762),
            .I(N__26755));
    LocalMux I__4323 (
            .O(N__26759),
            .I(N__26752));
    InMux I__4322 (
            .O(N__26758),
            .I(N__26749));
    LocalMux I__4321 (
            .O(N__26755),
            .I(N__26745));
    Span4Mux_h I__4320 (
            .O(N__26752),
            .I(N__26742));
    LocalMux I__4319 (
            .O(N__26749),
            .I(N__26739));
    InMux I__4318 (
            .O(N__26748),
            .I(N__26736));
    Span4Mux_v I__4317 (
            .O(N__26745),
            .I(N__26733));
    Span4Mux_v I__4316 (
            .O(N__26742),
            .I(N__26730));
    Span4Mux_h I__4315 (
            .O(N__26739),
            .I(N__26725));
    LocalMux I__4314 (
            .O(N__26736),
            .I(N__26725));
    Odrv4 I__4313 (
            .O(N__26733),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__4312 (
            .O(N__26730),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__4311 (
            .O(N__26725),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__4310 (
            .O(N__26718),
            .I(N__26713));
    InMux I__4309 (
            .O(N__26717),
            .I(N__26710));
    InMux I__4308 (
            .O(N__26716),
            .I(N__26707));
    LocalMux I__4307 (
            .O(N__26713),
            .I(N__26704));
    LocalMux I__4306 (
            .O(N__26710),
            .I(N__26701));
    LocalMux I__4305 (
            .O(N__26707),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    Odrv12 I__4304 (
            .O(N__26704),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    Odrv4 I__4303 (
            .O(N__26701),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    InMux I__4302 (
            .O(N__26694),
            .I(N__26688));
    InMux I__4301 (
            .O(N__26693),
            .I(N__26688));
    LocalMux I__4300 (
            .O(N__26688),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ));
    CascadeMux I__4299 (
            .O(N__26685),
            .I(N__26682));
    InMux I__4298 (
            .O(N__26682),
            .I(N__26679));
    LocalMux I__4297 (
            .O(N__26679),
            .I(N__26675));
    InMux I__4296 (
            .O(N__26678),
            .I(N__26672));
    Span4Mux_v I__4295 (
            .O(N__26675),
            .I(N__26669));
    LocalMux I__4294 (
            .O(N__26672),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    Odrv4 I__4293 (
            .O(N__26669),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    CascadeMux I__4292 (
            .O(N__26664),
            .I(N__26658));
    InMux I__4291 (
            .O(N__26663),
            .I(N__26653));
    InMux I__4290 (
            .O(N__26662),
            .I(N__26653));
    InMux I__4289 (
            .O(N__26661),
            .I(N__26650));
    InMux I__4288 (
            .O(N__26658),
            .I(N__26647));
    LocalMux I__4287 (
            .O(N__26653),
            .I(N__26644));
    LocalMux I__4286 (
            .O(N__26650),
            .I(N__26639));
    LocalMux I__4285 (
            .O(N__26647),
            .I(N__26639));
    Span4Mux_h I__4284 (
            .O(N__26644),
            .I(N__26636));
    Span4Mux_v I__4283 (
            .O(N__26639),
            .I(N__26633));
    Odrv4 I__4282 (
            .O(N__26636),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__4281 (
            .O(N__26633),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    CascadeMux I__4280 (
            .O(N__26628),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12_cascade_));
    InMux I__4279 (
            .O(N__26625),
            .I(N__26620));
    InMux I__4278 (
            .O(N__26624),
            .I(N__26617));
    InMux I__4277 (
            .O(N__26623),
            .I(N__26614));
    LocalMux I__4276 (
            .O(N__26620),
            .I(N__26611));
    LocalMux I__4275 (
            .O(N__26617),
            .I(N__26608));
    LocalMux I__4274 (
            .O(N__26614),
            .I(N__26603));
    Span4Mux_v I__4273 (
            .O(N__26611),
            .I(N__26603));
    Span4Mux_v I__4272 (
            .O(N__26608),
            .I(N__26600));
    Odrv4 I__4271 (
            .O(N__26603),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    Odrv4 I__4270 (
            .O(N__26600),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    InMux I__4269 (
            .O(N__26595),
            .I(N__26591));
    InMux I__4268 (
            .O(N__26594),
            .I(N__26587));
    LocalMux I__4267 (
            .O(N__26591),
            .I(N__26584));
    InMux I__4266 (
            .O(N__26590),
            .I(N__26581));
    LocalMux I__4265 (
            .O(N__26587),
            .I(N__26575));
    Span4Mux_v I__4264 (
            .O(N__26584),
            .I(N__26575));
    LocalMux I__4263 (
            .O(N__26581),
            .I(N__26572));
    InMux I__4262 (
            .O(N__26580),
            .I(N__26569));
    Span4Mux_h I__4261 (
            .O(N__26575),
            .I(N__26566));
    Span4Mux_v I__4260 (
            .O(N__26572),
            .I(N__26561));
    LocalMux I__4259 (
            .O(N__26569),
            .I(N__26561));
    Odrv4 I__4258 (
            .O(N__26566),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    Odrv4 I__4257 (
            .O(N__26561),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__4256 (
            .O(N__26556),
            .I(N__26550));
    InMux I__4255 (
            .O(N__26555),
            .I(N__26550));
    LocalMux I__4254 (
            .O(N__26550),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    InMux I__4253 (
            .O(N__26547),
            .I(N__26544));
    LocalMux I__4252 (
            .O(N__26544),
            .I(N__26540));
    InMux I__4251 (
            .O(N__26543),
            .I(N__26536));
    Span4Mux_v I__4250 (
            .O(N__26540),
            .I(N__26533));
    InMux I__4249 (
            .O(N__26539),
            .I(N__26530));
    LocalMux I__4248 (
            .O(N__26536),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    Odrv4 I__4247 (
            .O(N__26533),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    LocalMux I__4246 (
            .O(N__26530),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    CascadeMux I__4245 (
            .O(N__26523),
            .I(N__26518));
    InMux I__4244 (
            .O(N__26522),
            .I(N__26515));
    InMux I__4243 (
            .O(N__26521),
            .I(N__26511));
    InMux I__4242 (
            .O(N__26518),
            .I(N__26508));
    LocalMux I__4241 (
            .O(N__26515),
            .I(N__26505));
    InMux I__4240 (
            .O(N__26514),
            .I(N__26502));
    LocalMux I__4239 (
            .O(N__26511),
            .I(N__26499));
    LocalMux I__4238 (
            .O(N__26508),
            .I(N__26496));
    Span4Mux_h I__4237 (
            .O(N__26505),
            .I(N__26493));
    LocalMux I__4236 (
            .O(N__26502),
            .I(N__26490));
    Span4Mux_v I__4235 (
            .O(N__26499),
            .I(N__26487));
    Span4Mux_v I__4234 (
            .O(N__26496),
            .I(N__26484));
    Odrv4 I__4233 (
            .O(N__26493),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv12 I__4232 (
            .O(N__26490),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv4 I__4231 (
            .O(N__26487),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv4 I__4230 (
            .O(N__26484),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    CascadeMux I__4229 (
            .O(N__26475),
            .I(N__26472));
    InMux I__4228 (
            .O(N__26472),
            .I(N__26466));
    InMux I__4227 (
            .O(N__26471),
            .I(N__26466));
    LocalMux I__4226 (
            .O(N__26466),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    InMux I__4225 (
            .O(N__26463),
            .I(N__26460));
    LocalMux I__4224 (
            .O(N__26460),
            .I(N__26455));
    InMux I__4223 (
            .O(N__26459),
            .I(N__26452));
    InMux I__4222 (
            .O(N__26458),
            .I(N__26449));
    Span4Mux_h I__4221 (
            .O(N__26455),
            .I(N__26446));
    LocalMux I__4220 (
            .O(N__26452),
            .I(N__26443));
    LocalMux I__4219 (
            .O(N__26449),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    Odrv4 I__4218 (
            .O(N__26446),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    Odrv12 I__4217 (
            .O(N__26443),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    InMux I__4216 (
            .O(N__26436),
            .I(N__26432));
    InMux I__4215 (
            .O(N__26435),
            .I(N__26429));
    LocalMux I__4214 (
            .O(N__26432),
            .I(N__26426));
    LocalMux I__4213 (
            .O(N__26429),
            .I(N__26419));
    Span4Mux_v I__4212 (
            .O(N__26426),
            .I(N__26419));
    InMux I__4211 (
            .O(N__26425),
            .I(N__26414));
    InMux I__4210 (
            .O(N__26424),
            .I(N__26414));
    Span4Mux_v I__4209 (
            .O(N__26419),
            .I(N__26409));
    LocalMux I__4208 (
            .O(N__26414),
            .I(N__26409));
    Odrv4 I__4207 (
            .O(N__26409),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__4206 (
            .O(N__26406),
            .I(N__26402));
    InMux I__4205 (
            .O(N__26405),
            .I(N__26399));
    LocalMux I__4204 (
            .O(N__26402),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    LocalMux I__4203 (
            .O(N__26399),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    CascadeMux I__4202 (
            .O(N__26394),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11_cascade_));
    InMux I__4201 (
            .O(N__26391),
            .I(N__26383));
    InMux I__4200 (
            .O(N__26390),
            .I(N__26383));
    InMux I__4199 (
            .O(N__26389),
            .I(N__26378));
    InMux I__4198 (
            .O(N__26388),
            .I(N__26378));
    LocalMux I__4197 (
            .O(N__26383),
            .I(N__26375));
    LocalMux I__4196 (
            .O(N__26378),
            .I(N__26372));
    Span4Mux_v I__4195 (
            .O(N__26375),
            .I(N__26369));
    Odrv4 I__4194 (
            .O(N__26372),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    Odrv4 I__4193 (
            .O(N__26369),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__4192 (
            .O(N__26364),
            .I(N__26360));
    InMux I__4191 (
            .O(N__26363),
            .I(N__26357));
    LocalMux I__4190 (
            .O(N__26360),
            .I(N__26352));
    LocalMux I__4189 (
            .O(N__26357),
            .I(N__26349));
    InMux I__4188 (
            .O(N__26356),
            .I(N__26346));
    InMux I__4187 (
            .O(N__26355),
            .I(N__26343));
    Span4Mux_h I__4186 (
            .O(N__26352),
            .I(N__26340));
    Span4Mux_v I__4185 (
            .O(N__26349),
            .I(N__26335));
    LocalMux I__4184 (
            .O(N__26346),
            .I(N__26335));
    LocalMux I__4183 (
            .O(N__26343),
            .I(N__26332));
    Span4Mux_v I__4182 (
            .O(N__26340),
            .I(N__26327));
    Span4Mux_h I__4181 (
            .O(N__26335),
            .I(N__26327));
    Span4Mux_v I__4180 (
            .O(N__26332),
            .I(N__26324));
    Odrv4 I__4179 (
            .O(N__26327),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__4178 (
            .O(N__26324),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__4177 (
            .O(N__26319),
            .I(N__26316));
    LocalMux I__4176 (
            .O(N__26316),
            .I(N__26313));
    Span4Mux_h I__4175 (
            .O(N__26313),
            .I(N__26308));
    InMux I__4174 (
            .O(N__26312),
            .I(N__26305));
    InMux I__4173 (
            .O(N__26311),
            .I(N__26302));
    Span4Mux_v I__4172 (
            .O(N__26308),
            .I(N__26299));
    LocalMux I__4171 (
            .O(N__26305),
            .I(N__26296));
    LocalMux I__4170 (
            .O(N__26302),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__4169 (
            .O(N__26299),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__4168 (
            .O(N__26296),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    InMux I__4167 (
            .O(N__26289),
            .I(N__26283));
    InMux I__4166 (
            .O(N__26288),
            .I(N__26278));
    InMux I__4165 (
            .O(N__26287),
            .I(N__26278));
    InMux I__4164 (
            .O(N__26286),
            .I(N__26275));
    LocalMux I__4163 (
            .O(N__26283),
            .I(N__26272));
    LocalMux I__4162 (
            .O(N__26278),
            .I(N__26269));
    LocalMux I__4161 (
            .O(N__26275),
            .I(N__26266));
    Span4Mux_h I__4160 (
            .O(N__26272),
            .I(N__26261));
    Span4Mux_h I__4159 (
            .O(N__26269),
            .I(N__26261));
    Span4Mux_h I__4158 (
            .O(N__26266),
            .I(N__26258));
    Odrv4 I__4157 (
            .O(N__26261),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv4 I__4156 (
            .O(N__26258),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__4155 (
            .O(N__26253),
            .I(N__26247));
    InMux I__4154 (
            .O(N__26252),
            .I(N__26247));
    LocalMux I__4153 (
            .O(N__26247),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    InMux I__4152 (
            .O(N__26244),
            .I(N__26240));
    InMux I__4151 (
            .O(N__26243),
            .I(N__26236));
    LocalMux I__4150 (
            .O(N__26240),
            .I(N__26233));
    InMux I__4149 (
            .O(N__26239),
            .I(N__26230));
    LocalMux I__4148 (
            .O(N__26236),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    Odrv12 I__4147 (
            .O(N__26233),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__4146 (
            .O(N__26230),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    InMux I__4145 (
            .O(N__26223),
            .I(N__26219));
    InMux I__4144 (
            .O(N__26222),
            .I(N__26214));
    LocalMux I__4143 (
            .O(N__26219),
            .I(N__26211));
    InMux I__4142 (
            .O(N__26218),
            .I(N__26208));
    InMux I__4141 (
            .O(N__26217),
            .I(N__26205));
    LocalMux I__4140 (
            .O(N__26214),
            .I(N__26202));
    Span4Mux_v I__4139 (
            .O(N__26211),
            .I(N__26195));
    LocalMux I__4138 (
            .O(N__26208),
            .I(N__26195));
    LocalMux I__4137 (
            .O(N__26205),
            .I(N__26195));
    Span4Mux_h I__4136 (
            .O(N__26202),
            .I(N__26190));
    Span4Mux_h I__4135 (
            .O(N__26195),
            .I(N__26190));
    Odrv4 I__4134 (
            .O(N__26190),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__4133 (
            .O(N__26187),
            .I(N__26181));
    InMux I__4132 (
            .O(N__26186),
            .I(N__26181));
    LocalMux I__4131 (
            .O(N__26181),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__4130 (
            .O(N__26178),
            .I(N__26171));
    InMux I__4129 (
            .O(N__26177),
            .I(N__26171));
    InMux I__4128 (
            .O(N__26176),
            .I(N__26167));
    LocalMux I__4127 (
            .O(N__26171),
            .I(N__26164));
    InMux I__4126 (
            .O(N__26170),
            .I(N__26161));
    LocalMux I__4125 (
            .O(N__26167),
            .I(N__26156));
    Span4Mux_v I__4124 (
            .O(N__26164),
            .I(N__26156));
    LocalMux I__4123 (
            .O(N__26161),
            .I(N__26153));
    Span4Mux_v I__4122 (
            .O(N__26156),
            .I(N__26150));
    Span4Mux_h I__4121 (
            .O(N__26153),
            .I(N__26147));
    Odrv4 I__4120 (
            .O(N__26150),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__4119 (
            .O(N__26147),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__4118 (
            .O(N__26142),
            .I(N__26139));
    LocalMux I__4117 (
            .O(N__26139),
            .I(N__26135));
    InMux I__4116 (
            .O(N__26138),
            .I(N__26132));
    Odrv4 I__4115 (
            .O(N__26135),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    LocalMux I__4114 (
            .O(N__26132),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    CascadeMux I__4113 (
            .O(N__26127),
            .I(N__26124));
    InMux I__4112 (
            .O(N__26124),
            .I(N__26118));
    InMux I__4111 (
            .O(N__26123),
            .I(N__26118));
    LocalMux I__4110 (
            .O(N__26118),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__4109 (
            .O(N__26115),
            .I(N__26111));
    InMux I__4108 (
            .O(N__26114),
            .I(N__26108));
    LocalMux I__4107 (
            .O(N__26111),
            .I(N__26105));
    LocalMux I__4106 (
            .O(N__26108),
            .I(N__26098));
    Span4Mux_v I__4105 (
            .O(N__26105),
            .I(N__26098));
    InMux I__4104 (
            .O(N__26104),
            .I(N__26095));
    InMux I__4103 (
            .O(N__26103),
            .I(N__26092));
    Odrv4 I__4102 (
            .O(N__26098),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__4101 (
            .O(N__26095),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__4100 (
            .O(N__26092),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__4099 (
            .O(N__26085),
            .I(N__26082));
    LocalMux I__4098 (
            .O(N__26082),
            .I(N__26077));
    InMux I__4097 (
            .O(N__26081),
            .I(N__26074));
    InMux I__4096 (
            .O(N__26080),
            .I(N__26071));
    Span4Mux_h I__4095 (
            .O(N__26077),
            .I(N__26068));
    LocalMux I__4094 (
            .O(N__26074),
            .I(N__26065));
    LocalMux I__4093 (
            .O(N__26071),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__4092 (
            .O(N__26068),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv12 I__4091 (
            .O(N__26065),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__4090 (
            .O(N__26058),
            .I(N__26053));
    InMux I__4089 (
            .O(N__26057),
            .I(N__26050));
    InMux I__4088 (
            .O(N__26056),
            .I(N__26047));
    LocalMux I__4087 (
            .O(N__26053),
            .I(N__26043));
    LocalMux I__4086 (
            .O(N__26050),
            .I(N__26040));
    LocalMux I__4085 (
            .O(N__26047),
            .I(N__26037));
    InMux I__4084 (
            .O(N__26046),
            .I(N__26034));
    Span4Mux_v I__4083 (
            .O(N__26043),
            .I(N__26031));
    Span4Mux_v I__4082 (
            .O(N__26040),
            .I(N__26028));
    Span4Mux_h I__4081 (
            .O(N__26037),
            .I(N__26025));
    LocalMux I__4080 (
            .O(N__26034),
            .I(N__26022));
    Odrv4 I__4079 (
            .O(N__26031),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__4078 (
            .O(N__26028),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__4077 (
            .O(N__26025),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__4076 (
            .O(N__26022),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__4075 (
            .O(N__26013),
            .I(N__26009));
    InMux I__4074 (
            .O(N__26012),
            .I(N__26005));
    LocalMux I__4073 (
            .O(N__26009),
            .I(N__26002));
    InMux I__4072 (
            .O(N__26008),
            .I(N__25999));
    LocalMux I__4071 (
            .O(N__26005),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    Odrv4 I__4070 (
            .O(N__26002),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    LocalMux I__4069 (
            .O(N__25999),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    InMux I__4068 (
            .O(N__25992),
            .I(N__25989));
    LocalMux I__4067 (
            .O(N__25989),
            .I(N__25986));
    Odrv12 I__4066 (
            .O(N__25986),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ));
    InMux I__4065 (
            .O(N__25983),
            .I(N__25978));
    InMux I__4064 (
            .O(N__25982),
            .I(N__25974));
    InMux I__4063 (
            .O(N__25981),
            .I(N__25971));
    LocalMux I__4062 (
            .O(N__25978),
            .I(N__25968));
    InMux I__4061 (
            .O(N__25977),
            .I(N__25965));
    LocalMux I__4060 (
            .O(N__25974),
            .I(N__25962));
    LocalMux I__4059 (
            .O(N__25971),
            .I(N__25957));
    Span4Mux_h I__4058 (
            .O(N__25968),
            .I(N__25957));
    LocalMux I__4057 (
            .O(N__25965),
            .I(N__25954));
    Span4Mux_v I__4056 (
            .O(N__25962),
            .I(N__25947));
    Span4Mux_v I__4055 (
            .O(N__25957),
            .I(N__25947));
    Span4Mux_v I__4054 (
            .O(N__25954),
            .I(N__25947));
    Odrv4 I__4053 (
            .O(N__25947),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__4052 (
            .O(N__25944),
            .I(N__25941));
    LocalMux I__4051 (
            .O(N__25941),
            .I(N__25938));
    Odrv4 I__4050 (
            .O(N__25938),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ));
    InMux I__4049 (
            .O(N__25935),
            .I(N__25932));
    LocalMux I__4048 (
            .O(N__25932),
            .I(N__25929));
    Odrv4 I__4047 (
            .O(N__25929),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    CascadeMux I__4046 (
            .O(N__25926),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23_cascade_ ));
    InMux I__4045 (
            .O(N__25923),
            .I(N__25920));
    LocalMux I__4044 (
            .O(N__25920),
            .I(N__25917));
    Odrv4 I__4043 (
            .O(N__25917),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    CascadeMux I__4042 (
            .O(N__25914),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    InMux I__4041 (
            .O(N__25911),
            .I(N__25908));
    LocalMux I__4040 (
            .O(N__25908),
            .I(N__25903));
    InMux I__4039 (
            .O(N__25907),
            .I(N__25900));
    InMux I__4038 (
            .O(N__25906),
            .I(N__25897));
    Span4Mux_v I__4037 (
            .O(N__25903),
            .I(N__25894));
    LocalMux I__4036 (
            .O(N__25900),
            .I(N__25891));
    LocalMux I__4035 (
            .O(N__25897),
            .I(N__25886));
    Span4Mux_v I__4034 (
            .O(N__25894),
            .I(N__25886));
    Span4Mux_h I__4033 (
            .O(N__25891),
            .I(N__25883));
    Odrv4 I__4032 (
            .O(N__25886),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv4 I__4031 (
            .O(N__25883),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    InMux I__4030 (
            .O(N__25878),
            .I(N__25875));
    LocalMux I__4029 (
            .O(N__25875),
            .I(N__25871));
    InMux I__4028 (
            .O(N__25874),
            .I(N__25868));
    Span4Mux_v I__4027 (
            .O(N__25871),
            .I(N__25861));
    LocalMux I__4026 (
            .O(N__25868),
            .I(N__25861));
    InMux I__4025 (
            .O(N__25867),
            .I(N__25858));
    InMux I__4024 (
            .O(N__25866),
            .I(N__25855));
    Span4Mux_h I__4023 (
            .O(N__25861),
            .I(N__25850));
    LocalMux I__4022 (
            .O(N__25858),
            .I(N__25850));
    LocalMux I__4021 (
            .O(N__25855),
            .I(N__25847));
    Odrv4 I__4020 (
            .O(N__25850),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv4 I__4019 (
            .O(N__25847),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__4018 (
            .O(N__25842),
            .I(N__25836));
    InMux I__4017 (
            .O(N__25841),
            .I(N__25836));
    LocalMux I__4016 (
            .O(N__25836),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    InMux I__4015 (
            .O(N__25833),
            .I(N__25830));
    LocalMux I__4014 (
            .O(N__25830),
            .I(N__25827));
    Span4Mux_v I__4013 (
            .O(N__25827),
            .I(N__25823));
    InMux I__4012 (
            .O(N__25826),
            .I(N__25820));
    Odrv4 I__4011 (
            .O(N__25823),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__4010 (
            .O(N__25820),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    CascadeMux I__4009 (
            .O(N__25815),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_));
    InMux I__4008 (
            .O(N__25812),
            .I(N__25806));
    InMux I__4007 (
            .O(N__25811),
            .I(N__25806));
    LocalMux I__4006 (
            .O(N__25806),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ));
    InMux I__4005 (
            .O(N__25803),
            .I(N__25797));
    InMux I__4004 (
            .O(N__25802),
            .I(N__25797));
    LocalMux I__4003 (
            .O(N__25797),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ));
    InMux I__4002 (
            .O(N__25794),
            .I(N__25791));
    LocalMux I__4001 (
            .O(N__25791),
            .I(N__25788));
    Span4Mux_v I__4000 (
            .O(N__25788),
            .I(N__25783));
    InMux I__3999 (
            .O(N__25787),
            .I(N__25780));
    InMux I__3998 (
            .O(N__25786),
            .I(N__25777));
    Span4Mux_v I__3997 (
            .O(N__25783),
            .I(N__25772));
    LocalMux I__3996 (
            .O(N__25780),
            .I(N__25772));
    LocalMux I__3995 (
            .O(N__25777),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    Odrv4 I__3994 (
            .O(N__25772),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    CascadeMux I__3993 (
            .O(N__25767),
            .I(N__25763));
    InMux I__3992 (
            .O(N__25766),
            .I(N__25758));
    InMux I__3991 (
            .O(N__25763),
            .I(N__25758));
    LocalMux I__3990 (
            .O(N__25758),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    InMux I__3989 (
            .O(N__25755),
            .I(N__25749));
    InMux I__3988 (
            .O(N__25754),
            .I(N__25749));
    LocalMux I__3987 (
            .O(N__25749),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    CascadeMux I__3986 (
            .O(N__25746),
            .I(N__25742));
    InMux I__3985 (
            .O(N__25745),
            .I(N__25739));
    InMux I__3984 (
            .O(N__25742),
            .I(N__25736));
    LocalMux I__3983 (
            .O(N__25739),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    LocalMux I__3982 (
            .O(N__25736),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__3981 (
            .O(N__25731),
            .I(N__25727));
    InMux I__3980 (
            .O(N__25730),
            .I(N__25724));
    LocalMux I__3979 (
            .O(N__25727),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    LocalMux I__3978 (
            .O(N__25724),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__3977 (
            .O(N__25719),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__3976 (
            .O(N__25716),
            .I(N__25713));
    LocalMux I__3975 (
            .O(N__25713),
            .I(N__25709));
    InMux I__3974 (
            .O(N__25712),
            .I(N__25706));
    Odrv4 I__3973 (
            .O(N__25709),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    LocalMux I__3972 (
            .O(N__25706),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    CascadeMux I__3971 (
            .O(N__25701),
            .I(N__25696));
    InMux I__3970 (
            .O(N__25700),
            .I(N__25693));
    InMux I__3969 (
            .O(N__25699),
            .I(N__25690));
    InMux I__3968 (
            .O(N__25696),
            .I(N__25687));
    LocalMux I__3967 (
            .O(N__25693),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__3966 (
            .O(N__25690),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__3965 (
            .O(N__25687),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    InMux I__3964 (
            .O(N__25680),
            .I(N__25677));
    LocalMux I__3963 (
            .O(N__25677),
            .I(N__25674));
    Odrv4 I__3962 (
            .O(N__25674),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__3961 (
            .O(N__25671),
            .I(N__25665));
    InMux I__3960 (
            .O(N__25670),
            .I(N__25665));
    LocalMux I__3959 (
            .O(N__25665),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    CascadeMux I__3958 (
            .O(N__25662),
            .I(N__25659));
    InMux I__3957 (
            .O(N__25659),
            .I(N__25653));
    InMux I__3956 (
            .O(N__25658),
            .I(N__25653));
    LocalMux I__3955 (
            .O(N__25653),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    InMux I__3954 (
            .O(N__25650),
            .I(N__25646));
    InMux I__3953 (
            .O(N__25649),
            .I(N__25643));
    LocalMux I__3952 (
            .O(N__25646),
            .I(N__25640));
    LocalMux I__3951 (
            .O(N__25643),
            .I(N__25637));
    Span4Mux_v I__3950 (
            .O(N__25640),
            .I(N__25634));
    Span4Mux_h I__3949 (
            .O(N__25637),
            .I(N__25631));
    Span4Mux_h I__3948 (
            .O(N__25634),
            .I(N__25628));
    Span4Mux_h I__3947 (
            .O(N__25631),
            .I(N__25625));
    Span4Mux_h I__3946 (
            .O(N__25628),
            .I(N__25622));
    Odrv4 I__3945 (
            .O(N__25625),
            .I(\pwm_generator_inst.un3_threshold ));
    Odrv4 I__3944 (
            .O(N__25622),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__3943 (
            .O(N__25617),
            .I(N__25614));
    LocalMux I__3942 (
            .O(N__25614),
            .I(N__25611));
    Span4Mux_v I__3941 (
            .O(N__25611),
            .I(N__25608));
    Sp12to4 I__3940 (
            .O(N__25608),
            .I(N__25605));
    Odrv12 I__3939 (
            .O(N__25605),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__3938 (
            .O(N__25602),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__3937 (
            .O(N__25599),
            .I(N__25596));
    LocalMux I__3936 (
            .O(N__25596),
            .I(N__25593));
    Span4Mux_v I__3935 (
            .O(N__25593),
            .I(N__25590));
    Sp12to4 I__3934 (
            .O(N__25590),
            .I(N__25587));
    Odrv12 I__3933 (
            .O(N__25587),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__3932 (
            .O(N__25584),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__3931 (
            .O(N__25581),
            .I(N__25578));
    LocalMux I__3930 (
            .O(N__25578),
            .I(N__25575));
    Sp12to4 I__3929 (
            .O(N__25575),
            .I(N__25572));
    Span12Mux_s6_v I__3928 (
            .O(N__25572),
            .I(N__25569));
    Odrv12 I__3927 (
            .O(N__25569),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__3926 (
            .O(N__25566),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__3925 (
            .O(N__25563),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    InMux I__3924 (
            .O(N__25560),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__3923 (
            .O(N__25557),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__3922 (
            .O(N__25554),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__3921 (
            .O(N__25551),
            .I(bfn_9_27_0_));
    CEMux I__3920 (
            .O(N__25548),
            .I(N__25543));
    CEMux I__3919 (
            .O(N__25547),
            .I(N__25540));
    CEMux I__3918 (
            .O(N__25546),
            .I(N__25537));
    LocalMux I__3917 (
            .O(N__25543),
            .I(N__25533));
    LocalMux I__3916 (
            .O(N__25540),
            .I(N__25530));
    LocalMux I__3915 (
            .O(N__25537),
            .I(N__25527));
    CEMux I__3914 (
            .O(N__25536),
            .I(N__25524));
    Span4Mux_h I__3913 (
            .O(N__25533),
            .I(N__25521));
    Span4Mux_h I__3912 (
            .O(N__25530),
            .I(N__25518));
    Span4Mux_h I__3911 (
            .O(N__25527),
            .I(N__25515));
    LocalMux I__3910 (
            .O(N__25524),
            .I(N__25512));
    Odrv4 I__3909 (
            .O(N__25521),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    Odrv4 I__3908 (
            .O(N__25518),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    Odrv4 I__3907 (
            .O(N__25515),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    Odrv12 I__3906 (
            .O(N__25512),
            .I(\delay_measurement_inst.delay_hc_timer.N_199_i ));
    InMux I__3905 (
            .O(N__25503),
            .I(N__25500));
    LocalMux I__3904 (
            .O(N__25500),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__3903 (
            .O(N__25497),
            .I(N__25493));
    InMux I__3902 (
            .O(N__25496),
            .I(N__25490));
    LocalMux I__3901 (
            .O(N__25493),
            .I(\current_shift_inst.control_input_axb_0 ));
    LocalMux I__3900 (
            .O(N__25490),
            .I(\current_shift_inst.control_input_axb_0 ));
    InMux I__3899 (
            .O(N__25485),
            .I(N__25482));
    LocalMux I__3898 (
            .O(N__25482),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__3897 (
            .O(N__25479),
            .I(N__25476));
    LocalMux I__3896 (
            .O(N__25476),
            .I(\current_shift_inst.control_input_axb_3 ));
    CascadeMux I__3895 (
            .O(N__25473),
            .I(N__25468));
    InMux I__3894 (
            .O(N__25472),
            .I(N__25465));
    InMux I__3893 (
            .O(N__25471),
            .I(N__25462));
    InMux I__3892 (
            .O(N__25468),
            .I(N__25459));
    LocalMux I__3891 (
            .O(N__25465),
            .I(\current_shift_inst.N_1288_i ));
    LocalMux I__3890 (
            .O(N__25462),
            .I(\current_shift_inst.N_1288_i ));
    LocalMux I__3889 (
            .O(N__25459),
            .I(\current_shift_inst.N_1288_i ));
    InMux I__3888 (
            .O(N__25452),
            .I(N__25449));
    LocalMux I__3887 (
            .O(N__25449),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__3886 (
            .O(N__25446),
            .I(N__25443));
    LocalMux I__3885 (
            .O(N__25443),
            .I(\current_shift_inst.control_input_axb_7 ));
    CascadeMux I__3884 (
            .O(N__25440),
            .I(N__25437));
    InMux I__3883 (
            .O(N__25437),
            .I(N__25431));
    InMux I__3882 (
            .O(N__25436),
            .I(N__25431));
    LocalMux I__3881 (
            .O(N__25431),
            .I(N__25428));
    Odrv4 I__3880 (
            .O(N__25428),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ));
    InMux I__3879 (
            .O(N__25425),
            .I(N__25419));
    InMux I__3878 (
            .O(N__25424),
            .I(N__25419));
    LocalMux I__3877 (
            .O(N__25419),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ));
    InMux I__3876 (
            .O(N__25416),
            .I(N__25413));
    LocalMux I__3875 (
            .O(N__25413),
            .I(N__25410));
    Span4Mux_h I__3874 (
            .O(N__25410),
            .I(N__25406));
    InMux I__3873 (
            .O(N__25409),
            .I(N__25403));
    Odrv4 I__3872 (
            .O(N__25406),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    LocalMux I__3871 (
            .O(N__25403),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    CascadeMux I__3870 (
            .O(N__25398),
            .I(elapsed_time_ns_1_RNIK63T9_0_8_cascade_));
    InMux I__3869 (
            .O(N__25395),
            .I(N__25390));
    InMux I__3868 (
            .O(N__25394),
            .I(N__25385));
    InMux I__3867 (
            .O(N__25393),
            .I(N__25385));
    LocalMux I__3866 (
            .O(N__25390),
            .I(N__25381));
    LocalMux I__3865 (
            .O(N__25385),
            .I(N__25378));
    InMux I__3864 (
            .O(N__25384),
            .I(N__25375));
    Span4Mux_v I__3863 (
            .O(N__25381),
            .I(N__25370));
    Span4Mux_h I__3862 (
            .O(N__25378),
            .I(N__25370));
    LocalMux I__3861 (
            .O(N__25375),
            .I(N__25367));
    Odrv4 I__3860 (
            .O(N__25370),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__3859 (
            .O(N__25367),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__3858 (
            .O(N__25362),
            .I(N__25359));
    LocalMux I__3857 (
            .O(N__25359),
            .I(N__25356));
    Span12Mux_v I__3856 (
            .O(N__25356),
            .I(N__25353));
    Odrv12 I__3855 (
            .O(N__25353),
            .I(il_min_comp1_c));
    InMux I__3854 (
            .O(N__25350),
            .I(N__25338));
    InMux I__3853 (
            .O(N__25349),
            .I(N__25338));
    InMux I__3852 (
            .O(N__25348),
            .I(N__25338));
    InMux I__3851 (
            .O(N__25347),
            .I(N__25338));
    LocalMux I__3850 (
            .O(N__25338),
            .I(N__25309));
    InMux I__3849 (
            .O(N__25337),
            .I(N__25300));
    InMux I__3848 (
            .O(N__25336),
            .I(N__25300));
    InMux I__3847 (
            .O(N__25335),
            .I(N__25300));
    InMux I__3846 (
            .O(N__25334),
            .I(N__25300));
    InMux I__3845 (
            .O(N__25333),
            .I(N__25295));
    InMux I__3844 (
            .O(N__25332),
            .I(N__25295));
    InMux I__3843 (
            .O(N__25331),
            .I(N__25286));
    InMux I__3842 (
            .O(N__25330),
            .I(N__25286));
    InMux I__3841 (
            .O(N__25329),
            .I(N__25286));
    InMux I__3840 (
            .O(N__25328),
            .I(N__25286));
    InMux I__3839 (
            .O(N__25327),
            .I(N__25277));
    InMux I__3838 (
            .O(N__25326),
            .I(N__25277));
    InMux I__3837 (
            .O(N__25325),
            .I(N__25277));
    InMux I__3836 (
            .O(N__25324),
            .I(N__25277));
    InMux I__3835 (
            .O(N__25323),
            .I(N__25268));
    InMux I__3834 (
            .O(N__25322),
            .I(N__25268));
    InMux I__3833 (
            .O(N__25321),
            .I(N__25268));
    InMux I__3832 (
            .O(N__25320),
            .I(N__25268));
    InMux I__3831 (
            .O(N__25319),
            .I(N__25259));
    InMux I__3830 (
            .O(N__25318),
            .I(N__25259));
    InMux I__3829 (
            .O(N__25317),
            .I(N__25259));
    InMux I__3828 (
            .O(N__25316),
            .I(N__25259));
    InMux I__3827 (
            .O(N__25315),
            .I(N__25250));
    InMux I__3826 (
            .O(N__25314),
            .I(N__25250));
    InMux I__3825 (
            .O(N__25313),
            .I(N__25250));
    InMux I__3824 (
            .O(N__25312),
            .I(N__25250));
    Span4Mux_v I__3823 (
            .O(N__25309),
            .I(N__25247));
    LocalMux I__3822 (
            .O(N__25300),
            .I(N__25244));
    LocalMux I__3821 (
            .O(N__25295),
            .I(N__25241));
    LocalMux I__3820 (
            .O(N__25286),
            .I(N__25234));
    LocalMux I__3819 (
            .O(N__25277),
            .I(N__25234));
    LocalMux I__3818 (
            .O(N__25268),
            .I(N__25234));
    LocalMux I__3817 (
            .O(N__25259),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__3816 (
            .O(N__25250),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__3815 (
            .O(N__25247),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__3814 (
            .O(N__25244),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__3813 (
            .O(N__25241),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__3812 (
            .O(N__25234),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    CEMux I__3811 (
            .O(N__25221),
            .I(N__25214));
    CEMux I__3810 (
            .O(N__25220),
            .I(N__25211));
    CEMux I__3809 (
            .O(N__25219),
            .I(N__25208));
    CEMux I__3808 (
            .O(N__25218),
            .I(N__25205));
    CEMux I__3807 (
            .O(N__25217),
            .I(N__25202));
    LocalMux I__3806 (
            .O(N__25214),
            .I(N__25199));
    LocalMux I__3805 (
            .O(N__25211),
            .I(N__25196));
    LocalMux I__3804 (
            .O(N__25208),
            .I(N__25193));
    LocalMux I__3803 (
            .O(N__25205),
            .I(N__25190));
    LocalMux I__3802 (
            .O(N__25202),
            .I(N__25187));
    Span4Mux_h I__3801 (
            .O(N__25199),
            .I(N__25184));
    Span4Mux_v I__3800 (
            .O(N__25196),
            .I(N__25181));
    Span4Mux_v I__3799 (
            .O(N__25193),
            .I(N__25176));
    Span4Mux_h I__3798 (
            .O(N__25190),
            .I(N__25176));
    Span4Mux_h I__3797 (
            .O(N__25187),
            .I(N__25173));
    Odrv4 I__3796 (
            .O(N__25184),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    Odrv4 I__3795 (
            .O(N__25181),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    Odrv4 I__3794 (
            .O(N__25176),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    Odrv4 I__3793 (
            .O(N__25173),
            .I(\delay_measurement_inst.delay_hc_timer.N_198_i ));
    InMux I__3792 (
            .O(N__25164),
            .I(N__25160));
    InMux I__3791 (
            .O(N__25163),
            .I(N__25156));
    LocalMux I__3790 (
            .O(N__25160),
            .I(N__25153));
    InMux I__3789 (
            .O(N__25159),
            .I(N__25150));
    LocalMux I__3788 (
            .O(N__25156),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv4 I__3787 (
            .O(N__25153),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    LocalMux I__3786 (
            .O(N__25150),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    InMux I__3785 (
            .O(N__25143),
            .I(N__25140));
    LocalMux I__3784 (
            .O(N__25140),
            .I(N__25136));
    InMux I__3783 (
            .O(N__25139),
            .I(N__25133));
    Span4Mux_v I__3782 (
            .O(N__25136),
            .I(N__25128));
    LocalMux I__3781 (
            .O(N__25133),
            .I(N__25128));
    Span4Mux_v I__3780 (
            .O(N__25128),
            .I(N__25123));
    InMux I__3779 (
            .O(N__25127),
            .I(N__25120));
    InMux I__3778 (
            .O(N__25126),
            .I(N__25117));
    Odrv4 I__3777 (
            .O(N__25123),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__3776 (
            .O(N__25120),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__3775 (
            .O(N__25117),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__3774 (
            .O(N__25110),
            .I(N__25104));
    InMux I__3773 (
            .O(N__25109),
            .I(N__25104));
    LocalMux I__3772 (
            .O(N__25104),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    InMux I__3771 (
            .O(N__25101),
            .I(N__25097));
    InMux I__3770 (
            .O(N__25100),
            .I(N__25094));
    LocalMux I__3769 (
            .O(N__25097),
            .I(N__25090));
    LocalMux I__3768 (
            .O(N__25094),
            .I(N__25087));
    InMux I__3767 (
            .O(N__25093),
            .I(N__25084));
    Span4Mux_v I__3766 (
            .O(N__25090),
            .I(N__25081));
    Span4Mux_h I__3765 (
            .O(N__25087),
            .I(N__25078));
    LocalMux I__3764 (
            .O(N__25084),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    Odrv4 I__3763 (
            .O(N__25081),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    Odrv4 I__3762 (
            .O(N__25078),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    CascadeMux I__3761 (
            .O(N__25071),
            .I(N__25065));
    InMux I__3760 (
            .O(N__25070),
            .I(N__25062));
    InMux I__3759 (
            .O(N__25069),
            .I(N__25059));
    InMux I__3758 (
            .O(N__25068),
            .I(N__25056));
    InMux I__3757 (
            .O(N__25065),
            .I(N__25053));
    LocalMux I__3756 (
            .O(N__25062),
            .I(N__25050));
    LocalMux I__3755 (
            .O(N__25059),
            .I(N__25047));
    LocalMux I__3754 (
            .O(N__25056),
            .I(N__25042));
    LocalMux I__3753 (
            .O(N__25053),
            .I(N__25042));
    Span4Mux_h I__3752 (
            .O(N__25050),
            .I(N__25039));
    Span4Mux_h I__3751 (
            .O(N__25047),
            .I(N__25034));
    Span4Mux_h I__3750 (
            .O(N__25042),
            .I(N__25034));
    Odrv4 I__3749 (
            .O(N__25039),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__3748 (
            .O(N__25034),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    CascadeMux I__3747 (
            .O(N__25029),
            .I(N__25026));
    InMux I__3746 (
            .O(N__25026),
            .I(N__25020));
    InMux I__3745 (
            .O(N__25025),
            .I(N__25020));
    LocalMux I__3744 (
            .O(N__25020),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    InMux I__3743 (
            .O(N__25017),
            .I(N__25012));
    InMux I__3742 (
            .O(N__25016),
            .I(N__25006));
    InMux I__3741 (
            .O(N__25015),
            .I(N__25006));
    LocalMux I__3740 (
            .O(N__25012),
            .I(N__25003));
    InMux I__3739 (
            .O(N__25011),
            .I(N__25000));
    LocalMux I__3738 (
            .O(N__25006),
            .I(N__24997));
    Span4Mux_h I__3737 (
            .O(N__25003),
            .I(N__24992));
    LocalMux I__3736 (
            .O(N__25000),
            .I(N__24992));
    Odrv4 I__3735 (
            .O(N__24997),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__3734 (
            .O(N__24992),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__3733 (
            .O(N__24987),
            .I(N__24984));
    LocalMux I__3732 (
            .O(N__24984),
            .I(N__24981));
    Span4Mux_h I__3731 (
            .O(N__24981),
            .I(N__24977));
    InMux I__3730 (
            .O(N__24980),
            .I(N__24974));
    Odrv4 I__3729 (
            .O(N__24977),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__3728 (
            .O(N__24974),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    InMux I__3727 (
            .O(N__24969),
            .I(N__24966));
    LocalMux I__3726 (
            .O(N__24966),
            .I(N__24962));
    InMux I__3725 (
            .O(N__24965),
            .I(N__24958));
    Span4Mux_v I__3724 (
            .O(N__24962),
            .I(N__24955));
    InMux I__3723 (
            .O(N__24961),
            .I(N__24952));
    LocalMux I__3722 (
            .O(N__24958),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    Odrv4 I__3721 (
            .O(N__24955),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    LocalMux I__3720 (
            .O(N__24952),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    InMux I__3719 (
            .O(N__24945),
            .I(N__24941));
    CascadeMux I__3718 (
            .O(N__24944),
            .I(N__24936));
    LocalMux I__3717 (
            .O(N__24941),
            .I(N__24933));
    InMux I__3716 (
            .O(N__24940),
            .I(N__24930));
    InMux I__3715 (
            .O(N__24939),
            .I(N__24927));
    InMux I__3714 (
            .O(N__24936),
            .I(N__24924));
    Span4Mux_h I__3713 (
            .O(N__24933),
            .I(N__24921));
    LocalMux I__3712 (
            .O(N__24930),
            .I(N__24916));
    LocalMux I__3711 (
            .O(N__24927),
            .I(N__24916));
    LocalMux I__3710 (
            .O(N__24924),
            .I(N__24913));
    Odrv4 I__3709 (
            .O(N__24921),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__3708 (
            .O(N__24916),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__3707 (
            .O(N__24913),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__3706 (
            .O(N__24906),
            .I(N__24902));
    InMux I__3705 (
            .O(N__24905),
            .I(N__24898));
    LocalMux I__3704 (
            .O(N__24902),
            .I(N__24895));
    InMux I__3703 (
            .O(N__24901),
            .I(N__24892));
    LocalMux I__3702 (
            .O(N__24898),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    Odrv12 I__3701 (
            .O(N__24895),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    LocalMux I__3700 (
            .O(N__24892),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    InMux I__3699 (
            .O(N__24885),
            .I(N__24880));
    InMux I__3698 (
            .O(N__24884),
            .I(N__24877));
    InMux I__3697 (
            .O(N__24883),
            .I(N__24874));
    LocalMux I__3696 (
            .O(N__24880),
            .I(N__24870));
    LocalMux I__3695 (
            .O(N__24877),
            .I(N__24867));
    LocalMux I__3694 (
            .O(N__24874),
            .I(N__24864));
    InMux I__3693 (
            .O(N__24873),
            .I(N__24861));
    Span4Mux_v I__3692 (
            .O(N__24870),
            .I(N__24856));
    Span4Mux_v I__3691 (
            .O(N__24867),
            .I(N__24856));
    Span4Mux_h I__3690 (
            .O(N__24864),
            .I(N__24851));
    LocalMux I__3689 (
            .O(N__24861),
            .I(N__24851));
    Odrv4 I__3688 (
            .O(N__24856),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__3687 (
            .O(N__24851),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__3686 (
            .O(N__24846),
            .I(N__24843));
    LocalMux I__3685 (
            .O(N__24843),
            .I(N__24837));
    InMux I__3684 (
            .O(N__24842),
            .I(N__24834));
    InMux I__3683 (
            .O(N__24841),
            .I(N__24831));
    InMux I__3682 (
            .O(N__24840),
            .I(N__24828));
    Odrv4 I__3681 (
            .O(N__24837),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__3680 (
            .O(N__24834),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__3679 (
            .O(N__24831),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__3678 (
            .O(N__24828),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    InMux I__3677 (
            .O(N__24819),
            .I(N__24815));
    InMux I__3676 (
            .O(N__24818),
            .I(N__24811));
    LocalMux I__3675 (
            .O(N__24815),
            .I(N__24808));
    InMux I__3674 (
            .O(N__24814),
            .I(N__24805));
    LocalMux I__3673 (
            .O(N__24811),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__3672 (
            .O(N__24808),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    LocalMux I__3671 (
            .O(N__24805),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__3670 (
            .O(N__24798),
            .I(N__24794));
    InMux I__3669 (
            .O(N__24797),
            .I(N__24790));
    LocalMux I__3668 (
            .O(N__24794),
            .I(N__24787));
    InMux I__3667 (
            .O(N__24793),
            .I(N__24784));
    LocalMux I__3666 (
            .O(N__24790),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    Odrv12 I__3665 (
            .O(N__24787),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    LocalMux I__3664 (
            .O(N__24784),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    InMux I__3663 (
            .O(N__24777),
            .I(N__24773));
    InMux I__3662 (
            .O(N__24776),
            .I(N__24769));
    LocalMux I__3661 (
            .O(N__24773),
            .I(N__24765));
    InMux I__3660 (
            .O(N__24772),
            .I(N__24762));
    LocalMux I__3659 (
            .O(N__24769),
            .I(N__24759));
    InMux I__3658 (
            .O(N__24768),
            .I(N__24756));
    Span4Mux_h I__3657 (
            .O(N__24765),
            .I(N__24753));
    LocalMux I__3656 (
            .O(N__24762),
            .I(N__24750));
    Span4Mux_h I__3655 (
            .O(N__24759),
            .I(N__24747));
    LocalMux I__3654 (
            .O(N__24756),
            .I(N__24744));
    Span4Mux_v I__3653 (
            .O(N__24753),
            .I(N__24741));
    Span4Mux_h I__3652 (
            .O(N__24750),
            .I(N__24738));
    Span4Mux_v I__3651 (
            .O(N__24747),
            .I(N__24733));
    Span4Mux_h I__3650 (
            .O(N__24744),
            .I(N__24733));
    Odrv4 I__3649 (
            .O(N__24741),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__3648 (
            .O(N__24738),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__3647 (
            .O(N__24733),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__3646 (
            .O(N__24726),
            .I(N__24723));
    LocalMux I__3645 (
            .O(N__24723),
            .I(N__24719));
    InMux I__3644 (
            .O(N__24722),
            .I(N__24715));
    Span4Mux_v I__3643 (
            .O(N__24719),
            .I(N__24712));
    InMux I__3642 (
            .O(N__24718),
            .I(N__24709));
    LocalMux I__3641 (
            .O(N__24715),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    Odrv4 I__3640 (
            .O(N__24712),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    LocalMux I__3639 (
            .O(N__24709),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__3638 (
            .O(N__24702),
            .I(N__24698));
    InMux I__3637 (
            .O(N__24701),
            .I(N__24693));
    LocalMux I__3636 (
            .O(N__24698),
            .I(N__24690));
    InMux I__3635 (
            .O(N__24697),
            .I(N__24685));
    InMux I__3634 (
            .O(N__24696),
            .I(N__24685));
    LocalMux I__3633 (
            .O(N__24693),
            .I(N__24682));
    Span4Mux_h I__3632 (
            .O(N__24690),
            .I(N__24679));
    LocalMux I__3631 (
            .O(N__24685),
            .I(N__24676));
    Odrv4 I__3630 (
            .O(N__24682),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__3629 (
            .O(N__24679),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__3628 (
            .O(N__24676),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__3627 (
            .O(N__24669),
            .I(N__24665));
    InMux I__3626 (
            .O(N__24668),
            .I(N__24662));
    LocalMux I__3625 (
            .O(N__24665),
            .I(N__24657));
    LocalMux I__3624 (
            .O(N__24662),
            .I(N__24654));
    InMux I__3623 (
            .O(N__24661),
            .I(N__24649));
    InMux I__3622 (
            .O(N__24660),
            .I(N__24649));
    Span4Mux_v I__3621 (
            .O(N__24657),
            .I(N__24642));
    Span4Mux_v I__3620 (
            .O(N__24654),
            .I(N__24642));
    LocalMux I__3619 (
            .O(N__24649),
            .I(N__24642));
    Odrv4 I__3618 (
            .O(N__24642),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__3617 (
            .O(N__24639),
            .I(N__24634));
    InMux I__3616 (
            .O(N__24638),
            .I(N__24631));
    InMux I__3615 (
            .O(N__24637),
            .I(N__24628));
    LocalMux I__3614 (
            .O(N__24634),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    LocalMux I__3613 (
            .O(N__24631),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    LocalMux I__3612 (
            .O(N__24628),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    InMux I__3611 (
            .O(N__24621),
            .I(N__24617));
    InMux I__3610 (
            .O(N__24620),
            .I(N__24614));
    LocalMux I__3609 (
            .O(N__24617),
            .I(N__24609));
    LocalMux I__3608 (
            .O(N__24614),
            .I(N__24606));
    InMux I__3607 (
            .O(N__24613),
            .I(N__24601));
    InMux I__3606 (
            .O(N__24612),
            .I(N__24601));
    Span4Mux_v I__3605 (
            .O(N__24609),
            .I(N__24598));
    Span4Mux_h I__3604 (
            .O(N__24606),
            .I(N__24593));
    LocalMux I__3603 (
            .O(N__24601),
            .I(N__24593));
    Span4Mux_v I__3602 (
            .O(N__24598),
            .I(N__24590));
    Span4Mux_v I__3601 (
            .O(N__24593),
            .I(N__24587));
    Odrv4 I__3600 (
            .O(N__24590),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv4 I__3599 (
            .O(N__24587),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__3598 (
            .O(N__24582),
            .I(N__24578));
    InMux I__3597 (
            .O(N__24581),
            .I(N__24574));
    LocalMux I__3596 (
            .O(N__24578),
            .I(N__24571));
    InMux I__3595 (
            .O(N__24577),
            .I(N__24568));
    LocalMux I__3594 (
            .O(N__24574),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    Odrv4 I__3593 (
            .O(N__24571),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    LocalMux I__3592 (
            .O(N__24568),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    InMux I__3591 (
            .O(N__24561),
            .I(N__24557));
    InMux I__3590 (
            .O(N__24560),
            .I(N__24553));
    LocalMux I__3589 (
            .O(N__24557),
            .I(N__24550));
    InMux I__3588 (
            .O(N__24556),
            .I(N__24547));
    LocalMux I__3587 (
            .O(N__24553),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    Odrv4 I__3586 (
            .O(N__24550),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    LocalMux I__3585 (
            .O(N__24547),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    InMux I__3584 (
            .O(N__24540),
            .I(N__24537));
    LocalMux I__3583 (
            .O(N__24537),
            .I(N__24533));
    InMux I__3582 (
            .O(N__24536),
            .I(N__24530));
    Span4Mux_v I__3581 (
            .O(N__24533),
            .I(N__24526));
    LocalMux I__3580 (
            .O(N__24530),
            .I(N__24523));
    CascadeMux I__3579 (
            .O(N__24529),
            .I(N__24519));
    Span4Mux_h I__3578 (
            .O(N__24526),
            .I(N__24516));
    Span4Mux_h I__3577 (
            .O(N__24523),
            .I(N__24513));
    InMux I__3576 (
            .O(N__24522),
            .I(N__24508));
    InMux I__3575 (
            .O(N__24519),
            .I(N__24508));
    Odrv4 I__3574 (
            .O(N__24516),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__3573 (
            .O(N__24513),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    LocalMux I__3572 (
            .O(N__24508),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    CascadeMux I__3571 (
            .O(N__24501),
            .I(elapsed_time_ns_1_RNI68CN9_0_19_cascade_));
    CascadeMux I__3570 (
            .O(N__24498),
            .I(N__24495));
    InMux I__3569 (
            .O(N__24495),
            .I(N__24489));
    InMux I__3568 (
            .O(N__24494),
            .I(N__24489));
    LocalMux I__3567 (
            .O(N__24489),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__3566 (
            .O(N__24486),
            .I(N__24480));
    InMux I__3565 (
            .O(N__24485),
            .I(N__24480));
    LocalMux I__3564 (
            .O(N__24480),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    IoInMux I__3563 (
            .O(N__24477),
            .I(N__24474));
    LocalMux I__3562 (
            .O(N__24474),
            .I(GB_BUFFER_clock_output_0_THRU_CO));
    InMux I__3561 (
            .O(N__24471),
            .I(N__24468));
    LocalMux I__3560 (
            .O(N__24468),
            .I(N__24465));
    Glb2LocalMux I__3559 (
            .O(N__24465),
            .I(N__24462));
    GlobalMux I__3558 (
            .O(N__24462),
            .I(clk_12mhz));
    IoInMux I__3557 (
            .O(N__24459),
            .I(N__24456));
    LocalMux I__3556 (
            .O(N__24456),
            .I(N__24453));
    Span4Mux_s0_v I__3555 (
            .O(N__24453),
            .I(N__24450));
    Odrv4 I__3554 (
            .O(N__24450),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__3553 (
            .O(N__24447),
            .I(N__24444));
    LocalMux I__3552 (
            .O(N__24444),
            .I(N__24441));
    Odrv4 I__3551 (
            .O(N__24441),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__3550 (
            .O(N__24438),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__3549 (
            .O(N__24435),
            .I(N__24432));
    LocalMux I__3548 (
            .O(N__24432),
            .I(N__24429));
    Odrv4 I__3547 (
            .O(N__24429),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__3546 (
            .O(N__24426),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__3545 (
            .O(N__24423),
            .I(N__24420));
    LocalMux I__3544 (
            .O(N__24420),
            .I(N__24417));
    Odrv4 I__3543 (
            .O(N__24417),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__3542 (
            .O(N__24414),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__3541 (
            .O(N__24411),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__3540 (
            .O(N__24408),
            .I(N__24405));
    LocalMux I__3539 (
            .O(N__24405),
            .I(N__24401));
    InMux I__3538 (
            .O(N__24404),
            .I(N__24398));
    Odrv4 I__3537 (
            .O(N__24401),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__3536 (
            .O(N__24398),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__3535 (
            .O(N__24393),
            .I(N__24390));
    LocalMux I__3534 (
            .O(N__24390),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__3533 (
            .O(N__24387),
            .I(N__24384));
    LocalMux I__3532 (
            .O(N__24384),
            .I(N__24381));
    Span4Mux_h I__3531 (
            .O(N__24381),
            .I(N__24377));
    InMux I__3530 (
            .O(N__24380),
            .I(N__24374));
    Span4Mux_v I__3529 (
            .O(N__24377),
            .I(N__24371));
    LocalMux I__3528 (
            .O(N__24374),
            .I(N__24368));
    Span4Mux_h I__3527 (
            .O(N__24371),
            .I(N__24365));
    Odrv12 I__3526 (
            .O(N__24368),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv4 I__3525 (
            .O(N__24365),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    IoInMux I__3524 (
            .O(N__24360),
            .I(N__24357));
    LocalMux I__3523 (
            .O(N__24357),
            .I(N__24354));
    Span12Mux_s7_v I__3522 (
            .O(N__24354),
            .I(N__24351));
    Odrv12 I__3521 (
            .O(N__24351),
            .I(s4_phy_c));
    InMux I__3520 (
            .O(N__24348),
            .I(N__24345));
    LocalMux I__3519 (
            .O(N__24345),
            .I(N__24342));
    Odrv4 I__3518 (
            .O(N__24342),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__3517 (
            .O(N__24339),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__3516 (
            .O(N__24336),
            .I(N__24333));
    LocalMux I__3515 (
            .O(N__24333),
            .I(N__24330));
    Odrv4 I__3514 (
            .O(N__24330),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__3513 (
            .O(N__24327),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__3512 (
            .O(N__24324),
            .I(N__24321));
    LocalMux I__3511 (
            .O(N__24321),
            .I(N__24318));
    Odrv4 I__3510 (
            .O(N__24318),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__3509 (
            .O(N__24315),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__3508 (
            .O(N__24312),
            .I(N__24309));
    LocalMux I__3507 (
            .O(N__24309),
            .I(N__24306));
    Odrv4 I__3506 (
            .O(N__24306),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__3505 (
            .O(N__24303),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__3504 (
            .O(N__24300),
            .I(N__24297));
    LocalMux I__3503 (
            .O(N__24297),
            .I(N__24294));
    Odrv12 I__3502 (
            .O(N__24294),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__3501 (
            .O(N__24291),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__3500 (
            .O(N__24288),
            .I(N__24285));
    LocalMux I__3499 (
            .O(N__24285),
            .I(N__24282));
    Odrv12 I__3498 (
            .O(N__24282),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__3497 (
            .O(N__24279),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__3496 (
            .O(N__24276),
            .I(N__24273));
    LocalMux I__3495 (
            .O(N__24273),
            .I(N__24270));
    Odrv12 I__3494 (
            .O(N__24270),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__3493 (
            .O(N__24267),
            .I(bfn_8_16_0_));
    InMux I__3492 (
            .O(N__24264),
            .I(N__24261));
    LocalMux I__3491 (
            .O(N__24261),
            .I(N__24258));
    Odrv12 I__3490 (
            .O(N__24258),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__3489 (
            .O(N__24255),
            .I(\current_shift_inst.control_input_cry_8 ));
    CascadeMux I__3488 (
            .O(N__24252),
            .I(N__24248));
    CascadeMux I__3487 (
            .O(N__24251),
            .I(N__24245));
    InMux I__3486 (
            .O(N__24248),
            .I(N__24241));
    InMux I__3485 (
            .O(N__24245),
            .I(N__24238));
    InMux I__3484 (
            .O(N__24244),
            .I(N__24235));
    LocalMux I__3483 (
            .O(N__24241),
            .I(N__24232));
    LocalMux I__3482 (
            .O(N__24238),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__3481 (
            .O(N__24235),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__3480 (
            .O(N__24232),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__3479 (
            .O(N__24225),
            .I(bfn_8_14_0_));
    CascadeMux I__3478 (
            .O(N__24222),
            .I(N__24218));
    CascadeMux I__3477 (
            .O(N__24221),
            .I(N__24215));
    InMux I__3476 (
            .O(N__24218),
            .I(N__24211));
    InMux I__3475 (
            .O(N__24215),
            .I(N__24208));
    InMux I__3474 (
            .O(N__24214),
            .I(N__24205));
    LocalMux I__3473 (
            .O(N__24211),
            .I(N__24202));
    LocalMux I__3472 (
            .O(N__24208),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__3471 (
            .O(N__24205),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__3470 (
            .O(N__24202),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__3469 (
            .O(N__24195),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__3468 (
            .O(N__24192),
            .I(N__24189));
    InMux I__3467 (
            .O(N__24189),
            .I(N__24184));
    InMux I__3466 (
            .O(N__24188),
            .I(N__24181));
    InMux I__3465 (
            .O(N__24187),
            .I(N__24178));
    LocalMux I__3464 (
            .O(N__24184),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__3463 (
            .O(N__24181),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__3462 (
            .O(N__24178),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__3461 (
            .O(N__24171),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__3460 (
            .O(N__24168),
            .I(N__24165));
    InMux I__3459 (
            .O(N__24165),
            .I(N__24160));
    InMux I__3458 (
            .O(N__24164),
            .I(N__24157));
    InMux I__3457 (
            .O(N__24163),
            .I(N__24154));
    LocalMux I__3456 (
            .O(N__24160),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__3455 (
            .O(N__24157),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__3454 (
            .O(N__24154),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__3453 (
            .O(N__24147),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__3452 (
            .O(N__24144),
            .I(N__24140));
    InMux I__3451 (
            .O(N__24143),
            .I(N__24137));
    LocalMux I__3450 (
            .O(N__24140),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__3449 (
            .O(N__24137),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__3448 (
            .O(N__24132),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__3447 (
            .O(N__24129),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__3446 (
            .O(N__24126),
            .I(N__24122));
    InMux I__3445 (
            .O(N__24125),
            .I(N__24119));
    LocalMux I__3444 (
            .O(N__24122),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__3443 (
            .O(N__24119),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    InMux I__3442 (
            .O(N__24114),
            .I(N__24111));
    LocalMux I__3441 (
            .O(N__24111),
            .I(N__24108));
    Odrv12 I__3440 (
            .O(N__24108),
            .I(\current_shift_inst.control_input_18 ));
    InMux I__3439 (
            .O(N__24105),
            .I(N__24102));
    LocalMux I__3438 (
            .O(N__24102),
            .I(N__24099));
    Odrv12 I__3437 (
            .O(N__24099),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__3436 (
            .O(N__24096),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__3435 (
            .O(N__24093),
            .I(N__24088));
    InMux I__3434 (
            .O(N__24092),
            .I(N__24083));
    InMux I__3433 (
            .O(N__24091),
            .I(N__24083));
    LocalMux I__3432 (
            .O(N__24088),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__3431 (
            .O(N__24083),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__3430 (
            .O(N__24078),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__3429 (
            .O(N__24075),
            .I(N__24071));
    CascadeMux I__3428 (
            .O(N__24074),
            .I(N__24068));
    InMux I__3427 (
            .O(N__24071),
            .I(N__24064));
    InMux I__3426 (
            .O(N__24068),
            .I(N__24061));
    InMux I__3425 (
            .O(N__24067),
            .I(N__24058));
    LocalMux I__3424 (
            .O(N__24064),
            .I(N__24055));
    LocalMux I__3423 (
            .O(N__24061),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__3422 (
            .O(N__24058),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__3421 (
            .O(N__24055),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__3420 (
            .O(N__24048),
            .I(bfn_8_13_0_));
    CascadeMux I__3419 (
            .O(N__24045),
            .I(N__24041));
    CascadeMux I__3418 (
            .O(N__24044),
            .I(N__24038));
    InMux I__3417 (
            .O(N__24041),
            .I(N__24034));
    InMux I__3416 (
            .O(N__24038),
            .I(N__24031));
    InMux I__3415 (
            .O(N__24037),
            .I(N__24028));
    LocalMux I__3414 (
            .O(N__24034),
            .I(N__24025));
    LocalMux I__3413 (
            .O(N__24031),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__3412 (
            .O(N__24028),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__3411 (
            .O(N__24025),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__3410 (
            .O(N__24018),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__3409 (
            .O(N__24015),
            .I(N__24010));
    InMux I__3408 (
            .O(N__24014),
            .I(N__24005));
    InMux I__3407 (
            .O(N__24013),
            .I(N__24005));
    LocalMux I__3406 (
            .O(N__24010),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__3405 (
            .O(N__24005),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__3404 (
            .O(N__24000),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__3403 (
            .O(N__23997),
            .I(N__23994));
    InMux I__3402 (
            .O(N__23994),
            .I(N__23989));
    InMux I__3401 (
            .O(N__23993),
            .I(N__23986));
    InMux I__3400 (
            .O(N__23992),
            .I(N__23983));
    LocalMux I__3399 (
            .O(N__23989),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__3398 (
            .O(N__23986),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__3397 (
            .O(N__23983),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__3396 (
            .O(N__23976),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    CascadeMux I__3395 (
            .O(N__23973),
            .I(N__23968));
    CascadeMux I__3394 (
            .O(N__23972),
            .I(N__23965));
    InMux I__3393 (
            .O(N__23971),
            .I(N__23962));
    InMux I__3392 (
            .O(N__23968),
            .I(N__23957));
    InMux I__3391 (
            .O(N__23965),
            .I(N__23957));
    LocalMux I__3390 (
            .O(N__23962),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__3389 (
            .O(N__23957),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__3388 (
            .O(N__23952),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__3387 (
            .O(N__23949),
            .I(N__23946));
    InMux I__3386 (
            .O(N__23946),
            .I(N__23941));
    InMux I__3385 (
            .O(N__23945),
            .I(N__23938));
    InMux I__3384 (
            .O(N__23944),
            .I(N__23935));
    LocalMux I__3383 (
            .O(N__23941),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__3382 (
            .O(N__23938),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__3381 (
            .O(N__23935),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__3380 (
            .O(N__23928),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__3379 (
            .O(N__23925),
            .I(N__23920));
    InMux I__3378 (
            .O(N__23924),
            .I(N__23915));
    InMux I__3377 (
            .O(N__23923),
            .I(N__23915));
    LocalMux I__3376 (
            .O(N__23920),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__3375 (
            .O(N__23915),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__3374 (
            .O(N__23910),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__3373 (
            .O(N__23907),
            .I(N__23902));
    InMux I__3372 (
            .O(N__23906),
            .I(N__23897));
    InMux I__3371 (
            .O(N__23905),
            .I(N__23897));
    LocalMux I__3370 (
            .O(N__23902),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__3369 (
            .O(N__23897),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__3368 (
            .O(N__23892),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__3367 (
            .O(N__23889),
            .I(N__23884));
    InMux I__3366 (
            .O(N__23888),
            .I(N__23879));
    InMux I__3365 (
            .O(N__23887),
            .I(N__23879));
    LocalMux I__3364 (
            .O(N__23884),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__3363 (
            .O(N__23879),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__3362 (
            .O(N__23874),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__3361 (
            .O(N__23871),
            .I(N__23867));
    CascadeMux I__3360 (
            .O(N__23870),
            .I(N__23864));
    InMux I__3359 (
            .O(N__23867),
            .I(N__23860));
    InMux I__3358 (
            .O(N__23864),
            .I(N__23857));
    InMux I__3357 (
            .O(N__23863),
            .I(N__23854));
    LocalMux I__3356 (
            .O(N__23860),
            .I(N__23851));
    LocalMux I__3355 (
            .O(N__23857),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__3354 (
            .O(N__23854),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__3353 (
            .O(N__23851),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__3352 (
            .O(N__23844),
            .I(bfn_8_12_0_));
    CascadeMux I__3351 (
            .O(N__23841),
            .I(N__23837));
    CascadeMux I__3350 (
            .O(N__23840),
            .I(N__23834));
    InMux I__3349 (
            .O(N__23837),
            .I(N__23830));
    InMux I__3348 (
            .O(N__23834),
            .I(N__23827));
    InMux I__3347 (
            .O(N__23833),
            .I(N__23824));
    LocalMux I__3346 (
            .O(N__23830),
            .I(N__23821));
    LocalMux I__3345 (
            .O(N__23827),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__3344 (
            .O(N__23824),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__3343 (
            .O(N__23821),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__3342 (
            .O(N__23814),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__3341 (
            .O(N__23811),
            .I(N__23806));
    InMux I__3340 (
            .O(N__23810),
            .I(N__23801));
    InMux I__3339 (
            .O(N__23809),
            .I(N__23801));
    LocalMux I__3338 (
            .O(N__23806),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__3337 (
            .O(N__23801),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__3336 (
            .O(N__23796),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    CascadeMux I__3335 (
            .O(N__23793),
            .I(N__23790));
    InMux I__3334 (
            .O(N__23790),
            .I(N__23785));
    InMux I__3333 (
            .O(N__23789),
            .I(N__23782));
    InMux I__3332 (
            .O(N__23788),
            .I(N__23779));
    LocalMux I__3331 (
            .O(N__23785),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__3330 (
            .O(N__23782),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__3329 (
            .O(N__23779),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__3328 (
            .O(N__23772),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    CascadeMux I__3327 (
            .O(N__23769),
            .I(N__23764));
    CascadeMux I__3326 (
            .O(N__23768),
            .I(N__23761));
    InMux I__3325 (
            .O(N__23767),
            .I(N__23758));
    InMux I__3324 (
            .O(N__23764),
            .I(N__23753));
    InMux I__3323 (
            .O(N__23761),
            .I(N__23753));
    LocalMux I__3322 (
            .O(N__23758),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__3321 (
            .O(N__23753),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__3320 (
            .O(N__23748),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    CascadeMux I__3319 (
            .O(N__23745),
            .I(N__23742));
    InMux I__3318 (
            .O(N__23742),
            .I(N__23737));
    InMux I__3317 (
            .O(N__23741),
            .I(N__23734));
    InMux I__3316 (
            .O(N__23740),
            .I(N__23731));
    LocalMux I__3315 (
            .O(N__23737),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__3314 (
            .O(N__23734),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__3313 (
            .O(N__23731),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__3312 (
            .O(N__23724),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__3311 (
            .O(N__23721),
            .I(N__23716));
    InMux I__3310 (
            .O(N__23720),
            .I(N__23711));
    InMux I__3309 (
            .O(N__23719),
            .I(N__23711));
    LocalMux I__3308 (
            .O(N__23716),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__3307 (
            .O(N__23711),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__3306 (
            .O(N__23706),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    CascadeMux I__3305 (
            .O(N__23703),
            .I(N__23699));
    InMux I__3304 (
            .O(N__23702),
            .I(N__23695));
    InMux I__3303 (
            .O(N__23699),
            .I(N__23692));
    InMux I__3302 (
            .O(N__23698),
            .I(N__23689));
    LocalMux I__3301 (
            .O(N__23695),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__3300 (
            .O(N__23692),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__3299 (
            .O(N__23689),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__3298 (
            .O(N__23682),
            .I(bfn_8_11_0_));
    CascadeMux I__3297 (
            .O(N__23679),
            .I(N__23675));
    InMux I__3296 (
            .O(N__23678),
            .I(N__23671));
    InMux I__3295 (
            .O(N__23675),
            .I(N__23668));
    InMux I__3294 (
            .O(N__23674),
            .I(N__23665));
    LocalMux I__3293 (
            .O(N__23671),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__3292 (
            .O(N__23668),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__3291 (
            .O(N__23665),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__3290 (
            .O(N__23658),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__3289 (
            .O(N__23655),
            .I(N__23650));
    InMux I__3288 (
            .O(N__23654),
            .I(N__23645));
    InMux I__3287 (
            .O(N__23653),
            .I(N__23645));
    LocalMux I__3286 (
            .O(N__23650),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__3285 (
            .O(N__23645),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__3284 (
            .O(N__23640),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    CascadeMux I__3283 (
            .O(N__23637),
            .I(N__23634));
    InMux I__3282 (
            .O(N__23634),
            .I(N__23629));
    InMux I__3281 (
            .O(N__23633),
            .I(N__23626));
    InMux I__3280 (
            .O(N__23632),
            .I(N__23623));
    LocalMux I__3279 (
            .O(N__23629),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__3278 (
            .O(N__23626),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__3277 (
            .O(N__23623),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__3276 (
            .O(N__23616),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__3275 (
            .O(N__23613),
            .I(N__23608));
    CascadeMux I__3274 (
            .O(N__23612),
            .I(N__23605));
    InMux I__3273 (
            .O(N__23611),
            .I(N__23602));
    InMux I__3272 (
            .O(N__23608),
            .I(N__23597));
    InMux I__3271 (
            .O(N__23605),
            .I(N__23597));
    LocalMux I__3270 (
            .O(N__23602),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__3269 (
            .O(N__23597),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__3268 (
            .O(N__23592),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__3267 (
            .O(N__23589),
            .I(N__23586));
    InMux I__3266 (
            .O(N__23586),
            .I(N__23581));
    InMux I__3265 (
            .O(N__23585),
            .I(N__23578));
    InMux I__3264 (
            .O(N__23584),
            .I(N__23575));
    LocalMux I__3263 (
            .O(N__23581),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__3262 (
            .O(N__23578),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__3261 (
            .O(N__23575),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__3260 (
            .O(N__23568),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__3259 (
            .O(N__23565),
            .I(N__23560));
    InMux I__3258 (
            .O(N__23564),
            .I(N__23555));
    InMux I__3257 (
            .O(N__23563),
            .I(N__23555));
    LocalMux I__3256 (
            .O(N__23560),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__3255 (
            .O(N__23555),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__3254 (
            .O(N__23550),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__3253 (
            .O(N__23547),
            .I(N__23544));
    LocalMux I__3252 (
            .O(N__23544),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    InMux I__3251 (
            .O(N__23541),
            .I(N__23538));
    LocalMux I__3250 (
            .O(N__23538),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ));
    InMux I__3249 (
            .O(N__23535),
            .I(N__23532));
    LocalMux I__3248 (
            .O(N__23532),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ));
    InMux I__3247 (
            .O(N__23529),
            .I(N__23526));
    LocalMux I__3246 (
            .O(N__23526),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    InMux I__3245 (
            .O(N__23523),
            .I(N__23519));
    InMux I__3244 (
            .O(N__23522),
            .I(N__23516));
    LocalMux I__3243 (
            .O(N__23519),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    LocalMux I__3242 (
            .O(N__23516),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    InMux I__3241 (
            .O(N__23511),
            .I(N__23505));
    InMux I__3240 (
            .O(N__23510),
            .I(N__23505));
    LocalMux I__3239 (
            .O(N__23505),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ));
    CascadeMux I__3238 (
            .O(N__23502),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_ ));
    InMux I__3237 (
            .O(N__23499),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__3236 (
            .O(N__23496),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    InMux I__3235 (
            .O(N__23493),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    InMux I__3234 (
            .O(N__23490),
            .I(bfn_7_28_0_));
    InMux I__3233 (
            .O(N__23487),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__3232 (
            .O(N__23484),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__3231 (
            .O(N__23481),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__3230 (
            .O(N__23478),
            .I(N__23475));
    LocalMux I__3229 (
            .O(N__23475),
            .I(N__23472));
    Odrv12 I__3228 (
            .O(N__23472),
            .I(il_max_comp1_c));
    InMux I__3227 (
            .O(N__23469),
            .I(N__23466));
    LocalMux I__3226 (
            .O(N__23466),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    InMux I__3225 (
            .O(N__23463),
            .I(N__23460));
    LocalMux I__3224 (
            .O(N__23460),
            .I(N__23457));
    Span4Mux_h I__3223 (
            .O(N__23457),
            .I(N__23454));
    Span4Mux_h I__3222 (
            .O(N__23454),
            .I(N__23451));
    Odrv4 I__3221 (
            .O(N__23451),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__3220 (
            .O(N__23448),
            .I(N__23445));
    LocalMux I__3219 (
            .O(N__23445),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__3218 (
            .O(N__23442),
            .I(N__23439));
    LocalMux I__3217 (
            .O(N__23439),
            .I(N__23436));
    Span4Mux_h I__3216 (
            .O(N__23436),
            .I(N__23433));
    Span4Mux_h I__3215 (
            .O(N__23433),
            .I(N__23430));
    Odrv4 I__3214 (
            .O(N__23430),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__3213 (
            .O(N__23427),
            .I(N__23424));
    LocalMux I__3212 (
            .O(N__23424),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__3211 (
            .O(N__23421),
            .I(N__23418));
    LocalMux I__3210 (
            .O(N__23418),
            .I(N__23415));
    Span4Mux_v I__3209 (
            .O(N__23415),
            .I(N__23412));
    Span4Mux_h I__3208 (
            .O(N__23412),
            .I(N__23409));
    Odrv4 I__3207 (
            .O(N__23409),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__3206 (
            .O(N__23406),
            .I(N__23403));
    LocalMux I__3205 (
            .O(N__23403),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__3204 (
            .O(N__23400),
            .I(N__23397));
    LocalMux I__3203 (
            .O(N__23397),
            .I(N__23394));
    Span4Mux_v I__3202 (
            .O(N__23394),
            .I(N__23391));
    Span4Mux_h I__3201 (
            .O(N__23391),
            .I(N__23388));
    Odrv4 I__3200 (
            .O(N__23388),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__3199 (
            .O(N__23385),
            .I(N__23382));
    LocalMux I__3198 (
            .O(N__23382),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__3197 (
            .O(N__23379),
            .I(N__23376));
    LocalMux I__3196 (
            .O(N__23376),
            .I(N__23373));
    Span12Mux_s6_v I__3195 (
            .O(N__23373),
            .I(N__23370));
    Odrv12 I__3194 (
            .O(N__23370),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__3193 (
            .O(N__23367),
            .I(N__23364));
    LocalMux I__3192 (
            .O(N__23364),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__3191 (
            .O(N__23361),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    InMux I__3190 (
            .O(N__23358),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    InMux I__3189 (
            .O(N__23355),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__3188 (
            .O(N__23352),
            .I(N__23349));
    LocalMux I__3187 (
            .O(N__23349),
            .I(N__23346));
    Odrv4 I__3186 (
            .O(N__23346),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__3185 (
            .O(N__23343),
            .I(N__23340));
    LocalMux I__3184 (
            .O(N__23340),
            .I(N__23337));
    Span4Mux_v I__3183 (
            .O(N__23337),
            .I(N__23334));
    Span4Mux_h I__3182 (
            .O(N__23334),
            .I(N__23331));
    Odrv4 I__3181 (
            .O(N__23331),
            .I(\pwm_generator_inst.O_0 ));
    CascadeMux I__3180 (
            .O(N__23328),
            .I(N__23325));
    InMux I__3179 (
            .O(N__23325),
            .I(N__23322));
    LocalMux I__3178 (
            .O(N__23322),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__3177 (
            .O(N__23319),
            .I(N__23316));
    LocalMux I__3176 (
            .O(N__23316),
            .I(N__23313));
    Span12Mux_s7_v I__3175 (
            .O(N__23313),
            .I(N__23310));
    Odrv12 I__3174 (
            .O(N__23310),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__3173 (
            .O(N__23307),
            .I(N__23304));
    LocalMux I__3172 (
            .O(N__23304),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__3171 (
            .O(N__23301),
            .I(N__23298));
    LocalMux I__3170 (
            .O(N__23298),
            .I(N__23295));
    Span4Mux_h I__3169 (
            .O(N__23295),
            .I(N__23292));
    Span4Mux_h I__3168 (
            .O(N__23292),
            .I(N__23289));
    Odrv4 I__3167 (
            .O(N__23289),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__3166 (
            .O(N__23286),
            .I(N__23283));
    LocalMux I__3165 (
            .O(N__23283),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__3164 (
            .O(N__23280),
            .I(N__23277));
    LocalMux I__3163 (
            .O(N__23277),
            .I(N__23274));
    Span4Mux_h I__3162 (
            .O(N__23274),
            .I(N__23271));
    Span4Mux_h I__3161 (
            .O(N__23271),
            .I(N__23268));
    Odrv4 I__3160 (
            .O(N__23268),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__3159 (
            .O(N__23265),
            .I(N__23262));
    LocalMux I__3158 (
            .O(N__23262),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__3157 (
            .O(N__23259),
            .I(N__23256));
    LocalMux I__3156 (
            .O(N__23256),
            .I(N__23253));
    Span4Mux_h I__3155 (
            .O(N__23253),
            .I(N__23250));
    Span4Mux_h I__3154 (
            .O(N__23250),
            .I(N__23247));
    Odrv4 I__3153 (
            .O(N__23247),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__3152 (
            .O(N__23244),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__3151 (
            .O(N__23241),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__3150 (
            .O(N__23238),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__3149 (
            .O(N__23235),
            .I(bfn_7_13_0_));
    InMux I__3148 (
            .O(N__23232),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__3147 (
            .O(N__23229),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__3146 (
            .O(N__23226),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__3145 (
            .O(N__23223),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__3144 (
            .O(N__23220),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__3143 (
            .O(N__23217),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__3142 (
            .O(N__23214),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__3141 (
            .O(N__23211),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__3140 (
            .O(N__23208),
            .I(bfn_7_12_0_));
    InMux I__3139 (
            .O(N__23205),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__3138 (
            .O(N__23202),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__3137 (
            .O(N__23199),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__3136 (
            .O(N__23196),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__3135 (
            .O(N__23193),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__3134 (
            .O(N__23190),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__3133 (
            .O(N__23187),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__3132 (
            .O(N__23184),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__3131 (
            .O(N__23181),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__3130 (
            .O(N__23178),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__3129 (
            .O(N__23175),
            .I(bfn_7_11_0_));
    InMux I__3128 (
            .O(N__23172),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__3127 (
            .O(N__23169),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__3126 (
            .O(N__23166),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__3125 (
            .O(N__23163),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__3124 (
            .O(N__23160),
            .I(N__23128));
    InMux I__3123 (
            .O(N__23159),
            .I(N__23128));
    InMux I__3122 (
            .O(N__23158),
            .I(N__23128));
    InMux I__3121 (
            .O(N__23157),
            .I(N__23128));
    InMux I__3120 (
            .O(N__23156),
            .I(N__23128));
    InMux I__3119 (
            .O(N__23155),
            .I(N__23128));
    InMux I__3118 (
            .O(N__23154),
            .I(N__23128));
    InMux I__3117 (
            .O(N__23153),
            .I(N__23128));
    InMux I__3116 (
            .O(N__23152),
            .I(N__23111));
    InMux I__3115 (
            .O(N__23151),
            .I(N__23111));
    InMux I__3114 (
            .O(N__23150),
            .I(N__23111));
    InMux I__3113 (
            .O(N__23149),
            .I(N__23111));
    InMux I__3112 (
            .O(N__23148),
            .I(N__23111));
    InMux I__3111 (
            .O(N__23147),
            .I(N__23111));
    InMux I__3110 (
            .O(N__23146),
            .I(N__23111));
    InMux I__3109 (
            .O(N__23145),
            .I(N__23111));
    LocalMux I__3108 (
            .O(N__23128),
            .I(N__23107));
    LocalMux I__3107 (
            .O(N__23111),
            .I(N__23104));
    InMux I__3106 (
            .O(N__23110),
            .I(N__23101));
    Span4Mux_v I__3105 (
            .O(N__23107),
            .I(N__23098));
    Span4Mux_v I__3104 (
            .O(N__23104),
            .I(N__23095));
    LocalMux I__3103 (
            .O(N__23101),
            .I(N__23092));
    Span4Mux_v I__3102 (
            .O(N__23098),
            .I(N__23086));
    Span4Mux_v I__3101 (
            .O(N__23095),
            .I(N__23086));
    Span4Mux_s2_h I__3100 (
            .O(N__23092),
            .I(N__23083));
    InMux I__3099 (
            .O(N__23091),
            .I(N__23080));
    Span4Mux_h I__3098 (
            .O(N__23086),
            .I(N__23077));
    Span4Mux_v I__3097 (
            .O(N__23083),
            .I(N__23074));
    LocalMux I__3096 (
            .O(N__23080),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__3095 (
            .O(N__23077),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__3094 (
            .O(N__23074),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__3093 (
            .O(N__23067),
            .I(N__23063));
    InMux I__3092 (
            .O(N__23066),
            .I(N__23060));
    LocalMux I__3091 (
            .O(N__23063),
            .I(N__23057));
    LocalMux I__3090 (
            .O(N__23060),
            .I(N__23054));
    Span12Mux_v I__3089 (
            .O(N__23057),
            .I(N__23051));
    Odrv4 I__3088 (
            .O(N__23054),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv12 I__3087 (
            .O(N__23051),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__3086 (
            .O(N__23046),
            .I(N__23043));
    LocalMux I__3085 (
            .O(N__23043),
            .I(N__23040));
    Odrv12 I__3084 (
            .O(N__23040),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__3083 (
            .O(N__23037),
            .I(elapsed_time_ns_1_RNI02CN9_0_13_cascade_));
    InMux I__3082 (
            .O(N__23034),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__3081 (
            .O(N__23031),
            .I(N__23028));
    LocalMux I__3080 (
            .O(N__23028),
            .I(N__23024));
    InMux I__3079 (
            .O(N__23027),
            .I(N__23021));
    Span4Mux_s1_h I__3078 (
            .O(N__23024),
            .I(N__23018));
    LocalMux I__3077 (
            .O(N__23021),
            .I(N__23015));
    Span4Mux_h I__3076 (
            .O(N__23018),
            .I(N__23012));
    Odrv4 I__3075 (
            .O(N__23015),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__3074 (
            .O(N__23012),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__3073 (
            .O(N__23007),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__3072 (
            .O(N__23004),
            .I(N__23000));
    InMux I__3071 (
            .O(N__23003),
            .I(N__22997));
    LocalMux I__3070 (
            .O(N__23000),
            .I(N__22994));
    LocalMux I__3069 (
            .O(N__22997),
            .I(N__22991));
    Span4Mux_s1_h I__3068 (
            .O(N__22994),
            .I(N__22988));
    Span4Mux_h I__3067 (
            .O(N__22991),
            .I(N__22983));
    Span4Mux_h I__3066 (
            .O(N__22988),
            .I(N__22983));
    Odrv4 I__3065 (
            .O(N__22983),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__3064 (
            .O(N__22980),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__3063 (
            .O(N__22977),
            .I(N__22974));
    LocalMux I__3062 (
            .O(N__22974),
            .I(N__22970));
    InMux I__3061 (
            .O(N__22973),
            .I(N__22967));
    Span12Mux_s5_h I__3060 (
            .O(N__22970),
            .I(N__22964));
    LocalMux I__3059 (
            .O(N__22967),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv12 I__3058 (
            .O(N__22964),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__3057 (
            .O(N__22959),
            .I(bfn_5_16_0_));
    InMux I__3056 (
            .O(N__22956),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__3055 (
            .O(N__22953),
            .I(N__22950));
    LocalMux I__3054 (
            .O(N__22950),
            .I(N__22946));
    InMux I__3053 (
            .O(N__22949),
            .I(N__22943));
    Span4Mux_s1_h I__3052 (
            .O(N__22946),
            .I(N__22940));
    LocalMux I__3051 (
            .O(N__22943),
            .I(N__22937));
    Span4Mux_h I__3050 (
            .O(N__22940),
            .I(N__22934));
    Odrv4 I__3049 (
            .O(N__22937),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__3048 (
            .O(N__22934),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__3047 (
            .O(N__22929),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__3046 (
            .O(N__22926),
            .I(N__22923));
    LocalMux I__3045 (
            .O(N__22923),
            .I(N__22919));
    InMux I__3044 (
            .O(N__22922),
            .I(N__22916));
    Span4Mux_s1_h I__3043 (
            .O(N__22919),
            .I(N__22913));
    LocalMux I__3042 (
            .O(N__22916),
            .I(N__22910));
    Span4Mux_h I__3041 (
            .O(N__22913),
            .I(N__22907));
    Odrv4 I__3040 (
            .O(N__22910),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__3039 (
            .O(N__22907),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__3038 (
            .O(N__22902),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__3037 (
            .O(N__22899),
            .I(N__22896));
    LocalMux I__3036 (
            .O(N__22896),
            .I(N__22893));
    Span4Mux_s1_h I__3035 (
            .O(N__22893),
            .I(N__22889));
    InMux I__3034 (
            .O(N__22892),
            .I(N__22886));
    Span4Mux_h I__3033 (
            .O(N__22889),
            .I(N__22883));
    LocalMux I__3032 (
            .O(N__22886),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__3031 (
            .O(N__22883),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__3030 (
            .O(N__22878),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__3029 (
            .O(N__22875),
            .I(N__22872));
    LocalMux I__3028 (
            .O(N__22872),
            .I(N__22868));
    InMux I__3027 (
            .O(N__22871),
            .I(N__22865));
    Span4Mux_s1_h I__3026 (
            .O(N__22868),
            .I(N__22862));
    LocalMux I__3025 (
            .O(N__22865),
            .I(N__22859));
    Span4Mux_h I__3024 (
            .O(N__22862),
            .I(N__22856));
    Odrv4 I__3023 (
            .O(N__22859),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv4 I__3022 (
            .O(N__22856),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__3021 (
            .O(N__22851),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__3020 (
            .O(N__22848),
            .I(N__22845));
    LocalMux I__3019 (
            .O(N__22845),
            .I(N__22842));
    Odrv4 I__3018 (
            .O(N__22842),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__3017 (
            .O(N__22839),
            .I(N__22836));
    LocalMux I__3016 (
            .O(N__22836),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__3015 (
            .O(N__22833),
            .I(N__22828));
    InMux I__3014 (
            .O(N__22832),
            .I(N__22825));
    InMux I__3013 (
            .O(N__22831),
            .I(N__22822));
    LocalMux I__3012 (
            .O(N__22828),
            .I(N__22819));
    LocalMux I__3011 (
            .O(N__22825),
            .I(N__22816));
    LocalMux I__3010 (
            .O(N__22822),
            .I(N__22812));
    Span4Mux_v I__3009 (
            .O(N__22819),
            .I(N__22809));
    Span4Mux_v I__3008 (
            .O(N__22816),
            .I(N__22806));
    InMux I__3007 (
            .O(N__22815),
            .I(N__22803));
    Span4Mux_v I__3006 (
            .O(N__22812),
            .I(N__22800));
    Odrv4 I__3005 (
            .O(N__22809),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__3004 (
            .O(N__22806),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__3003 (
            .O(N__22803),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__3002 (
            .O(N__22800),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__3001 (
            .O(N__22791),
            .I(N__22787));
    InMux I__3000 (
            .O(N__22790),
            .I(N__22783));
    LocalMux I__2999 (
            .O(N__22787),
            .I(N__22780));
    InMux I__2998 (
            .O(N__22786),
            .I(N__22777));
    LocalMux I__2997 (
            .O(N__22783),
            .I(N__22774));
    Span4Mux_h I__2996 (
            .O(N__22780),
            .I(N__22768));
    LocalMux I__2995 (
            .O(N__22777),
            .I(N__22768));
    Span4Mux_h I__2994 (
            .O(N__22774),
            .I(N__22765));
    InMux I__2993 (
            .O(N__22773),
            .I(N__22762));
    Span4Mux_v I__2992 (
            .O(N__22768),
            .I(N__22759));
    Odrv4 I__2991 (
            .O(N__22765),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__2990 (
            .O(N__22762),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__2989 (
            .O(N__22759),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__2988 (
            .O(N__22752),
            .I(N__22748));
    CascadeMux I__2987 (
            .O(N__22751),
            .I(N__22745));
    InMux I__2986 (
            .O(N__22748),
            .I(N__22741));
    InMux I__2985 (
            .O(N__22745),
            .I(N__22738));
    InMux I__2984 (
            .O(N__22744),
            .I(N__22734));
    LocalMux I__2983 (
            .O(N__22741),
            .I(N__22731));
    LocalMux I__2982 (
            .O(N__22738),
            .I(N__22728));
    InMux I__2981 (
            .O(N__22737),
            .I(N__22725));
    LocalMux I__2980 (
            .O(N__22734),
            .I(N__22722));
    Span4Mux_h I__2979 (
            .O(N__22731),
            .I(N__22719));
    Span4Mux_h I__2978 (
            .O(N__22728),
            .I(N__22714));
    LocalMux I__2977 (
            .O(N__22725),
            .I(N__22714));
    Odrv4 I__2976 (
            .O(N__22722),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__2975 (
            .O(N__22719),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__2974 (
            .O(N__22714),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__2973 (
            .O(N__22707),
            .I(N__22688));
    InMux I__2972 (
            .O(N__22706),
            .I(N__22685));
    InMux I__2971 (
            .O(N__22705),
            .I(N__22682));
    InMux I__2970 (
            .O(N__22704),
            .I(N__22679));
    InMux I__2969 (
            .O(N__22703),
            .I(N__22668));
    InMux I__2968 (
            .O(N__22702),
            .I(N__22668));
    InMux I__2967 (
            .O(N__22701),
            .I(N__22668));
    InMux I__2966 (
            .O(N__22700),
            .I(N__22668));
    InMux I__2965 (
            .O(N__22699),
            .I(N__22668));
    InMux I__2964 (
            .O(N__22698),
            .I(N__22665));
    InMux I__2963 (
            .O(N__22697),
            .I(N__22661));
    InMux I__2962 (
            .O(N__22696),
            .I(N__22635));
    InMux I__2961 (
            .O(N__22695),
            .I(N__22635));
    InMux I__2960 (
            .O(N__22694),
            .I(N__22635));
    InMux I__2959 (
            .O(N__22693),
            .I(N__22635));
    InMux I__2958 (
            .O(N__22692),
            .I(N__22635));
    InMux I__2957 (
            .O(N__22691),
            .I(N__22635));
    LocalMux I__2956 (
            .O(N__22688),
            .I(N__22632));
    LocalMux I__2955 (
            .O(N__22685),
            .I(N__22621));
    LocalMux I__2954 (
            .O(N__22682),
            .I(N__22621));
    LocalMux I__2953 (
            .O(N__22679),
            .I(N__22621));
    LocalMux I__2952 (
            .O(N__22668),
            .I(N__22621));
    LocalMux I__2951 (
            .O(N__22665),
            .I(N__22621));
    InMux I__2950 (
            .O(N__22664),
            .I(N__22617));
    LocalMux I__2949 (
            .O(N__22661),
            .I(N__22614));
    InMux I__2948 (
            .O(N__22660),
            .I(N__22599));
    InMux I__2947 (
            .O(N__22659),
            .I(N__22599));
    InMux I__2946 (
            .O(N__22658),
            .I(N__22599));
    InMux I__2945 (
            .O(N__22657),
            .I(N__22599));
    InMux I__2944 (
            .O(N__22656),
            .I(N__22599));
    InMux I__2943 (
            .O(N__22655),
            .I(N__22599));
    InMux I__2942 (
            .O(N__22654),
            .I(N__22599));
    InMux I__2941 (
            .O(N__22653),
            .I(N__22596));
    InMux I__2940 (
            .O(N__22652),
            .I(N__22585));
    InMux I__2939 (
            .O(N__22651),
            .I(N__22585));
    InMux I__2938 (
            .O(N__22650),
            .I(N__22585));
    InMux I__2937 (
            .O(N__22649),
            .I(N__22585));
    InMux I__2936 (
            .O(N__22648),
            .I(N__22585));
    LocalMux I__2935 (
            .O(N__22635),
            .I(N__22582));
    Span4Mux_v I__2934 (
            .O(N__22632),
            .I(N__22577));
    Span4Mux_v I__2933 (
            .O(N__22621),
            .I(N__22577));
    InMux I__2932 (
            .O(N__22620),
            .I(N__22574));
    LocalMux I__2931 (
            .O(N__22617),
            .I(N__22569));
    Span4Mux_h I__2930 (
            .O(N__22614),
            .I(N__22569));
    LocalMux I__2929 (
            .O(N__22599),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__2928 (
            .O(N__22596),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__2927 (
            .O(N__22585),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__2926 (
            .O(N__22582),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__2925 (
            .O(N__22577),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__2924 (
            .O(N__22574),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__2923 (
            .O(N__22569),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__2922 (
            .O(N__22554),
            .I(N__22551));
    LocalMux I__2921 (
            .O(N__22551),
            .I(N__22548));
    Odrv12 I__2920 (
            .O(N__22548),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__2919 (
            .O(N__22545),
            .I(N__22542));
    LocalMux I__2918 (
            .O(N__22542),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__2917 (
            .O(N__22539),
            .I(N__22535));
    InMux I__2916 (
            .O(N__22538),
            .I(N__22532));
    LocalMux I__2915 (
            .O(N__22535),
            .I(N__22529));
    LocalMux I__2914 (
            .O(N__22532),
            .I(N__22524));
    Span12Mux_v I__2913 (
            .O(N__22529),
            .I(N__22524));
    Odrv12 I__2912 (
            .O(N__22524),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__2911 (
            .O(N__22521),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__2910 (
            .O(N__22518),
            .I(N__22515));
    LocalMux I__2909 (
            .O(N__22515),
            .I(N__22512));
    Span4Mux_s1_h I__2908 (
            .O(N__22512),
            .I(N__22508));
    InMux I__2907 (
            .O(N__22511),
            .I(N__22505));
    Span4Mux_h I__2906 (
            .O(N__22508),
            .I(N__22502));
    LocalMux I__2905 (
            .O(N__22505),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv4 I__2904 (
            .O(N__22502),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__2903 (
            .O(N__22497),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__2902 (
            .O(N__22494),
            .I(N__22491));
    LocalMux I__2901 (
            .O(N__22491),
            .I(N__22487));
    InMux I__2900 (
            .O(N__22490),
            .I(N__22484));
    Span4Mux_s1_h I__2899 (
            .O(N__22487),
            .I(N__22481));
    LocalMux I__2898 (
            .O(N__22484),
            .I(N__22478));
    Span4Mux_h I__2897 (
            .O(N__22481),
            .I(N__22475));
    Odrv4 I__2896 (
            .O(N__22478),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv4 I__2895 (
            .O(N__22475),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__2894 (
            .O(N__22470),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__2893 (
            .O(N__22467),
            .I(N__22463));
    InMux I__2892 (
            .O(N__22466),
            .I(N__22460));
    LocalMux I__2891 (
            .O(N__22463),
            .I(N__22457));
    LocalMux I__2890 (
            .O(N__22460),
            .I(N__22454));
    Span4Mux_v I__2889 (
            .O(N__22457),
            .I(N__22451));
    Span4Mux_v I__2888 (
            .O(N__22454),
            .I(N__22448));
    Sp12to4 I__2887 (
            .O(N__22451),
            .I(N__22445));
    Span4Mux_h I__2886 (
            .O(N__22448),
            .I(N__22442));
    Odrv12 I__2885 (
            .O(N__22445),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv4 I__2884 (
            .O(N__22442),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__2883 (
            .O(N__22437),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__2882 (
            .O(N__22434),
            .I(N__22430));
    InMux I__2881 (
            .O(N__22433),
            .I(N__22427));
    LocalMux I__2880 (
            .O(N__22430),
            .I(N__22424));
    LocalMux I__2879 (
            .O(N__22427),
            .I(N__22421));
    Span4Mux_v I__2878 (
            .O(N__22424),
            .I(N__22418));
    Span4Mux_v I__2877 (
            .O(N__22421),
            .I(N__22415));
    Span4Mux_h I__2876 (
            .O(N__22418),
            .I(N__22412));
    Odrv4 I__2875 (
            .O(N__22415),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv4 I__2874 (
            .O(N__22412),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__2873 (
            .O(N__22407),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__2872 (
            .O(N__22404),
            .I(N__22400));
    InMux I__2871 (
            .O(N__22403),
            .I(N__22397));
    LocalMux I__2870 (
            .O(N__22400),
            .I(N__22392));
    LocalMux I__2869 (
            .O(N__22397),
            .I(N__22392));
    Odrv4 I__2868 (
            .O(N__22392),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2867 (
            .O(N__22389),
            .I(N__22385));
    InMux I__2866 (
            .O(N__22388),
            .I(N__22382));
    LocalMux I__2865 (
            .O(N__22385),
            .I(N__22379));
    LocalMux I__2864 (
            .O(N__22382),
            .I(N__22376));
    Odrv4 I__2863 (
            .O(N__22379),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    Odrv4 I__2862 (
            .O(N__22376),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2861 (
            .O(N__22371),
            .I(N__22368));
    LocalMux I__2860 (
            .O(N__22368),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__2859 (
            .O(N__22365),
            .I(N__22361));
    InMux I__2858 (
            .O(N__22364),
            .I(N__22356));
    InMux I__2857 (
            .O(N__22361),
            .I(N__22356));
    LocalMux I__2856 (
            .O(N__22356),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2855 (
            .O(N__22353),
            .I(N__22347));
    InMux I__2854 (
            .O(N__22352),
            .I(N__22347));
    LocalMux I__2853 (
            .O(N__22347),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2852 (
            .O(N__22344),
            .I(N__22340));
    CascadeMux I__2851 (
            .O(N__22343),
            .I(N__22337));
    LocalMux I__2850 (
            .O(N__22340),
            .I(N__22334));
    InMux I__2849 (
            .O(N__22337),
            .I(N__22331));
    Odrv4 I__2848 (
            .O(N__22334),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__2847 (
            .O(N__22331),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2846 (
            .O(N__22326),
            .I(N__22322));
    InMux I__2845 (
            .O(N__22325),
            .I(N__22319));
    LocalMux I__2844 (
            .O(N__22322),
            .I(N__22316));
    LocalMux I__2843 (
            .O(N__22319),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    Odrv4 I__2842 (
            .O(N__22316),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    CascadeMux I__2841 (
            .O(N__22311),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ));
    InMux I__2840 (
            .O(N__22308),
            .I(N__22305));
    LocalMux I__2839 (
            .O(N__22305),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2838 (
            .O(N__22302),
            .I(N__22296));
    InMux I__2837 (
            .O(N__22301),
            .I(N__22296));
    LocalMux I__2836 (
            .O(N__22296),
            .I(N__22293));
    Odrv4 I__2835 (
            .O(N__22293),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2834 (
            .O(N__22290),
            .I(N__22284));
    InMux I__2833 (
            .O(N__22289),
            .I(N__22284));
    LocalMux I__2832 (
            .O(N__22284),
            .I(N__22281));
    Odrv4 I__2831 (
            .O(N__22281),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2830 (
            .O(N__22278),
            .I(N__22272));
    InMux I__2829 (
            .O(N__22277),
            .I(N__22272));
    LocalMux I__2828 (
            .O(N__22272),
            .I(N__22269));
    Odrv12 I__2827 (
            .O(N__22269),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    CascadeMux I__2826 (
            .O(N__22266),
            .I(N__22263));
    InMux I__2825 (
            .O(N__22263),
            .I(N__22257));
    InMux I__2824 (
            .O(N__22262),
            .I(N__22257));
    LocalMux I__2823 (
            .O(N__22257),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    CascadeMux I__2822 (
            .O(N__22254),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    InMux I__2821 (
            .O(N__22251),
            .I(N__22245));
    InMux I__2820 (
            .O(N__22250),
            .I(N__22245));
    LocalMux I__2819 (
            .O(N__22245),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2818 (
            .O(N__22242),
            .I(N__22239));
    LocalMux I__2817 (
            .O(N__22239),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__2816 (
            .O(N__22236),
            .I(N__22233));
    LocalMux I__2815 (
            .O(N__22233),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__2814 (
            .O(N__22230),
            .I(N__22219));
    CascadeMux I__2813 (
            .O(N__22229),
            .I(N__22215));
    CascadeMux I__2812 (
            .O(N__22228),
            .I(N__22211));
    CascadeMux I__2811 (
            .O(N__22227),
            .I(N__22208));
    CascadeMux I__2810 (
            .O(N__22226),
            .I(N__22204));
    CascadeMux I__2809 (
            .O(N__22225),
            .I(N__22200));
    CascadeMux I__2808 (
            .O(N__22224),
            .I(N__22196));
    InMux I__2807 (
            .O(N__22223),
            .I(N__22178));
    InMux I__2806 (
            .O(N__22222),
            .I(N__22178));
    InMux I__2805 (
            .O(N__22219),
            .I(N__22178));
    InMux I__2804 (
            .O(N__22218),
            .I(N__22178));
    InMux I__2803 (
            .O(N__22215),
            .I(N__22178));
    InMux I__2802 (
            .O(N__22214),
            .I(N__22178));
    InMux I__2801 (
            .O(N__22211),
            .I(N__22178));
    InMux I__2800 (
            .O(N__22208),
            .I(N__22161));
    InMux I__2799 (
            .O(N__22207),
            .I(N__22161));
    InMux I__2798 (
            .O(N__22204),
            .I(N__22161));
    InMux I__2797 (
            .O(N__22203),
            .I(N__22161));
    InMux I__2796 (
            .O(N__22200),
            .I(N__22161));
    InMux I__2795 (
            .O(N__22199),
            .I(N__22161));
    InMux I__2794 (
            .O(N__22196),
            .I(N__22161));
    InMux I__2793 (
            .O(N__22195),
            .I(N__22161));
    CascadeMux I__2792 (
            .O(N__22194),
            .I(N__22158));
    CascadeMux I__2791 (
            .O(N__22193),
            .I(N__22154));
    LocalMux I__2790 (
            .O(N__22178),
            .I(N__22149));
    LocalMux I__2789 (
            .O(N__22161),
            .I(N__22149));
    InMux I__2788 (
            .O(N__22158),
            .I(N__22142));
    InMux I__2787 (
            .O(N__22157),
            .I(N__22142));
    InMux I__2786 (
            .O(N__22154),
            .I(N__22142));
    Span4Mux_v I__2785 (
            .O(N__22149),
            .I(N__22137));
    LocalMux I__2784 (
            .O(N__22142),
            .I(N__22137));
    Odrv4 I__2783 (
            .O(N__22137),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__2782 (
            .O(N__22134),
            .I(N__22131));
    InMux I__2781 (
            .O(N__22131),
            .I(N__22128));
    LocalMux I__2780 (
            .O(N__22128),
            .I(N__22125));
    Odrv4 I__2779 (
            .O(N__22125),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__2778 (
            .O(N__22122),
            .I(N__22118));
    InMux I__2777 (
            .O(N__22121),
            .I(N__22114));
    LocalMux I__2776 (
            .O(N__22118),
            .I(N__22111));
    InMux I__2775 (
            .O(N__22117),
            .I(N__22107));
    LocalMux I__2774 (
            .O(N__22114),
            .I(N__22104));
    Span4Mux_v I__2773 (
            .O(N__22111),
            .I(N__22101));
    InMux I__2772 (
            .O(N__22110),
            .I(N__22098));
    LocalMux I__2771 (
            .O(N__22107),
            .I(N__22095));
    Span4Mux_v I__2770 (
            .O(N__22104),
            .I(N__22092));
    Odrv4 I__2769 (
            .O(N__22101),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__2768 (
            .O(N__22098),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__2767 (
            .O(N__22095),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__2766 (
            .O(N__22092),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__2765 (
            .O(N__22083),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    CascadeMux I__2764 (
            .O(N__22080),
            .I(N__22077));
    InMux I__2763 (
            .O(N__22077),
            .I(N__22073));
    InMux I__2762 (
            .O(N__22076),
            .I(N__22068));
    LocalMux I__2761 (
            .O(N__22073),
            .I(N__22065));
    InMux I__2760 (
            .O(N__22072),
            .I(N__22062));
    InMux I__2759 (
            .O(N__22071),
            .I(N__22059));
    LocalMux I__2758 (
            .O(N__22068),
            .I(N__22056));
    Span4Mux_v I__2757 (
            .O(N__22065),
            .I(N__22053));
    LocalMux I__2756 (
            .O(N__22062),
            .I(N__22050));
    LocalMux I__2755 (
            .O(N__22059),
            .I(N__22045));
    Span4Mux_v I__2754 (
            .O(N__22056),
            .I(N__22045));
    Odrv4 I__2753 (
            .O(N__22053),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv12 I__2752 (
            .O(N__22050),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__2751 (
            .O(N__22045),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__2750 (
            .O(N__22038),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2749 (
            .O(N__22035),
            .I(N__22031));
    InMux I__2748 (
            .O(N__22034),
            .I(N__22027));
    LocalMux I__2747 (
            .O(N__22031),
            .I(N__22023));
    CascadeMux I__2746 (
            .O(N__22030),
            .I(N__22020));
    LocalMux I__2745 (
            .O(N__22027),
            .I(N__22017));
    InMux I__2744 (
            .O(N__22026),
            .I(N__22014));
    Span4Mux_v I__2743 (
            .O(N__22023),
            .I(N__22011));
    InMux I__2742 (
            .O(N__22020),
            .I(N__22008));
    Sp12to4 I__2741 (
            .O(N__22017),
            .I(N__22003));
    LocalMux I__2740 (
            .O(N__22014),
            .I(N__22003));
    Odrv4 I__2739 (
            .O(N__22011),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__2738 (
            .O(N__22008),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv12 I__2737 (
            .O(N__22003),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__2736 (
            .O(N__21996),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    CascadeMux I__2735 (
            .O(N__21993),
            .I(N__21990));
    InMux I__2734 (
            .O(N__21990),
            .I(N__21987));
    LocalMux I__2733 (
            .O(N__21987),
            .I(N__21983));
    InMux I__2732 (
            .O(N__21986),
            .I(N__21978));
    Span4Mux_v I__2731 (
            .O(N__21983),
            .I(N__21975));
    InMux I__2730 (
            .O(N__21982),
            .I(N__21972));
    InMux I__2729 (
            .O(N__21981),
            .I(N__21969));
    LocalMux I__2728 (
            .O(N__21978),
            .I(N__21966));
    Odrv4 I__2727 (
            .O(N__21975),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__2726 (
            .O(N__21972),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__2725 (
            .O(N__21969),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__2724 (
            .O(N__21966),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__2723 (
            .O(N__21957),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2722 (
            .O(N__21954),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2721 (
            .O(N__21951),
            .I(N__21948));
    LocalMux I__2720 (
            .O(N__21948),
            .I(N__21945));
    Span4Mux_s3_h I__2719 (
            .O(N__21945),
            .I(N__21942));
    Odrv4 I__2718 (
            .O(N__21942),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2717 (
            .O(N__21939),
            .I(N__21936));
    LocalMux I__2716 (
            .O(N__21936),
            .I(N__21932));
    InMux I__2715 (
            .O(N__21935),
            .I(N__21929));
    Odrv4 I__2714 (
            .O(N__21932),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    LocalMux I__2713 (
            .O(N__21929),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2712 (
            .O(N__21924),
            .I(N__21921));
    LocalMux I__2711 (
            .O(N__21921),
            .I(N__21917));
    InMux I__2710 (
            .O(N__21920),
            .I(N__21914));
    Odrv4 I__2709 (
            .O(N__21917),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    LocalMux I__2708 (
            .O(N__21914),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2707 (
            .O(N__21909),
            .I(N__21906));
    LocalMux I__2706 (
            .O(N__21906),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__2705 (
            .O(N__21903),
            .I(N__21899));
    InMux I__2704 (
            .O(N__21902),
            .I(N__21896));
    LocalMux I__2703 (
            .O(N__21899),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__2702 (
            .O(N__21896),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    CascadeMux I__2701 (
            .O(N__21891),
            .I(N__21888));
    InMux I__2700 (
            .O(N__21888),
            .I(N__21884));
    InMux I__2699 (
            .O(N__21887),
            .I(N__21881));
    LocalMux I__2698 (
            .O(N__21884),
            .I(N__21878));
    LocalMux I__2697 (
            .O(N__21881),
            .I(N__21875));
    Odrv12 I__2696 (
            .O(N__21878),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    Odrv4 I__2695 (
            .O(N__21875),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2694 (
            .O(N__21870),
            .I(N__21867));
    LocalMux I__2693 (
            .O(N__21867),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__2692 (
            .O(N__21864),
            .I(N__21861));
    LocalMux I__2691 (
            .O(N__21861),
            .I(N__21855));
    CascadeMux I__2690 (
            .O(N__21860),
            .I(N__21852));
    InMux I__2689 (
            .O(N__21859),
            .I(N__21849));
    InMux I__2688 (
            .O(N__21858),
            .I(N__21846));
    Span4Mux_v I__2687 (
            .O(N__21855),
            .I(N__21843));
    InMux I__2686 (
            .O(N__21852),
            .I(N__21840));
    LocalMux I__2685 (
            .O(N__21849),
            .I(N__21835));
    LocalMux I__2684 (
            .O(N__21846),
            .I(N__21835));
    Odrv4 I__2683 (
            .O(N__21843),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__2682 (
            .O(N__21840),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__2681 (
            .O(N__21835),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__2680 (
            .O(N__21828),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    CascadeMux I__2679 (
            .O(N__21825),
            .I(N__21821));
    CascadeMux I__2678 (
            .O(N__21824),
            .I(N__21818));
    InMux I__2677 (
            .O(N__21821),
            .I(N__21814));
    InMux I__2676 (
            .O(N__21818),
            .I(N__21811));
    InMux I__2675 (
            .O(N__21817),
            .I(N__21808));
    LocalMux I__2674 (
            .O(N__21814),
            .I(N__21805));
    LocalMux I__2673 (
            .O(N__21811),
            .I(N__21799));
    LocalMux I__2672 (
            .O(N__21808),
            .I(N__21799));
    Span4Mux_v I__2671 (
            .O(N__21805),
            .I(N__21796));
    InMux I__2670 (
            .O(N__21804),
            .I(N__21793));
    Span4Mux_v I__2669 (
            .O(N__21799),
            .I(N__21790));
    Odrv4 I__2668 (
            .O(N__21796),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__2667 (
            .O(N__21793),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__2666 (
            .O(N__21790),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__2665 (
            .O(N__21783),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2664 (
            .O(N__21780),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__2663 (
            .O(N__21777),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2662 (
            .O(N__21774),
            .I(N__21770));
    InMux I__2661 (
            .O(N__21773),
            .I(N__21765));
    LocalMux I__2660 (
            .O(N__21770),
            .I(N__21762));
    InMux I__2659 (
            .O(N__21769),
            .I(N__21759));
    InMux I__2658 (
            .O(N__21768),
            .I(N__21756));
    LocalMux I__2657 (
            .O(N__21765),
            .I(N__21753));
    Span4Mux_v I__2656 (
            .O(N__21762),
            .I(N__21750));
    LocalMux I__2655 (
            .O(N__21759),
            .I(N__21747));
    LocalMux I__2654 (
            .O(N__21756),
            .I(N__21742));
    Span4Mux_v I__2653 (
            .O(N__21753),
            .I(N__21742));
    Odrv4 I__2652 (
            .O(N__21750),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv12 I__2651 (
            .O(N__21747),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__2650 (
            .O(N__21742),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__2649 (
            .O(N__21735),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    CascadeMux I__2648 (
            .O(N__21732),
            .I(N__21728));
    InMux I__2647 (
            .O(N__21731),
            .I(N__21725));
    InMux I__2646 (
            .O(N__21728),
            .I(N__21721));
    LocalMux I__2645 (
            .O(N__21725),
            .I(N__21717));
    InMux I__2644 (
            .O(N__21724),
            .I(N__21714));
    LocalMux I__2643 (
            .O(N__21721),
            .I(N__21711));
    CascadeMux I__2642 (
            .O(N__21720),
            .I(N__21708));
    Span4Mux_h I__2641 (
            .O(N__21717),
            .I(N__21703));
    LocalMux I__2640 (
            .O(N__21714),
            .I(N__21703));
    Span4Mux_v I__2639 (
            .O(N__21711),
            .I(N__21700));
    InMux I__2638 (
            .O(N__21708),
            .I(N__21697));
    Span4Mux_v I__2637 (
            .O(N__21703),
            .I(N__21694));
    Odrv4 I__2636 (
            .O(N__21700),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__2635 (
            .O(N__21697),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__2634 (
            .O(N__21694),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__2633 (
            .O(N__21687),
            .I(N__21684));
    InMux I__2632 (
            .O(N__21684),
            .I(N__21680));
    InMux I__2631 (
            .O(N__21683),
            .I(N__21677));
    LocalMux I__2630 (
            .O(N__21680),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    LocalMux I__2629 (
            .O(N__21677),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2628 (
            .O(N__21672),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2627 (
            .O(N__21669),
            .I(N__21665));
    InMux I__2626 (
            .O(N__21668),
            .I(N__21662));
    LocalMux I__2625 (
            .O(N__21665),
            .I(N__21659));
    LocalMux I__2624 (
            .O(N__21662),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    Odrv4 I__2623 (
            .O(N__21659),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2622 (
            .O(N__21654),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    CascadeMux I__2621 (
            .O(N__21651),
            .I(N__21647));
    InMux I__2620 (
            .O(N__21650),
            .I(N__21644));
    InMux I__2619 (
            .O(N__21647),
            .I(N__21640));
    LocalMux I__2618 (
            .O(N__21644),
            .I(N__21636));
    InMux I__2617 (
            .O(N__21643),
            .I(N__21633));
    LocalMux I__2616 (
            .O(N__21640),
            .I(N__21630));
    InMux I__2615 (
            .O(N__21639),
            .I(N__21627));
    Span4Mux_v I__2614 (
            .O(N__21636),
            .I(N__21622));
    LocalMux I__2613 (
            .O(N__21633),
            .I(N__21622));
    Span4Mux_v I__2612 (
            .O(N__21630),
            .I(N__21619));
    LocalMux I__2611 (
            .O(N__21627),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__2610 (
            .O(N__21622),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__2609 (
            .O(N__21619),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__2608 (
            .O(N__21612),
            .I(bfn_3_20_0_));
    CascadeMux I__2607 (
            .O(N__21609),
            .I(N__21605));
    CascadeMux I__2606 (
            .O(N__21608),
            .I(N__21602));
    InMux I__2605 (
            .O(N__21605),
            .I(N__21599));
    InMux I__2604 (
            .O(N__21602),
            .I(N__21596));
    LocalMux I__2603 (
            .O(N__21599),
            .I(N__21593));
    LocalMux I__2602 (
            .O(N__21596),
            .I(N__21588));
    Span4Mux_h I__2601 (
            .O(N__21593),
            .I(N__21585));
    InMux I__2600 (
            .O(N__21592),
            .I(N__21582));
    InMux I__2599 (
            .O(N__21591),
            .I(N__21579));
    Span4Mux_v I__2598 (
            .O(N__21588),
            .I(N__21576));
    Sp12to4 I__2597 (
            .O(N__21585),
            .I(N__21571));
    LocalMux I__2596 (
            .O(N__21582),
            .I(N__21571));
    LocalMux I__2595 (
            .O(N__21579),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__2594 (
            .O(N__21576),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv12 I__2593 (
            .O(N__21571),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__2592 (
            .O(N__21564),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2591 (
            .O(N__21561),
            .I(N__21558));
    LocalMux I__2590 (
            .O(N__21558),
            .I(N__21555));
    Odrv12 I__2589 (
            .O(N__21555),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__2588 (
            .O(N__21552),
            .I(N__21548));
    CascadeMux I__2587 (
            .O(N__21551),
            .I(N__21545));
    InMux I__2586 (
            .O(N__21548),
            .I(N__21542));
    InMux I__2585 (
            .O(N__21545),
            .I(N__21539));
    LocalMux I__2584 (
            .O(N__21542),
            .I(N__21536));
    LocalMux I__2583 (
            .O(N__21539),
            .I(N__21530));
    Span4Mux_h I__2582 (
            .O(N__21536),
            .I(N__21530));
    InMux I__2581 (
            .O(N__21535),
            .I(N__21526));
    Span4Mux_v I__2580 (
            .O(N__21530),
            .I(N__21523));
    InMux I__2579 (
            .O(N__21529),
            .I(N__21520));
    LocalMux I__2578 (
            .O(N__21526),
            .I(N__21517));
    Odrv4 I__2577 (
            .O(N__21523),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__2576 (
            .O(N__21520),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv12 I__2575 (
            .O(N__21517),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__2574 (
            .O(N__21510),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2573 (
            .O(N__21507),
            .I(N__21504));
    LocalMux I__2572 (
            .O(N__21504),
            .I(N__21501));
    Odrv4 I__2571 (
            .O(N__21501),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__2570 (
            .O(N__21498),
            .I(N__21495));
    InMux I__2569 (
            .O(N__21495),
            .I(N__21491));
    InMux I__2568 (
            .O(N__21494),
            .I(N__21488));
    LocalMux I__2567 (
            .O(N__21491),
            .I(N__21484));
    LocalMux I__2566 (
            .O(N__21488),
            .I(N__21481));
    InMux I__2565 (
            .O(N__21487),
            .I(N__21478));
    Span4Mux_v I__2564 (
            .O(N__21484),
            .I(N__21474));
    Span12Mux_s2_h I__2563 (
            .O(N__21481),
            .I(N__21469));
    LocalMux I__2562 (
            .O(N__21478),
            .I(N__21469));
    InMux I__2561 (
            .O(N__21477),
            .I(N__21466));
    Odrv4 I__2560 (
            .O(N__21474),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv12 I__2559 (
            .O(N__21469),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__2558 (
            .O(N__21466),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__2557 (
            .O(N__21459),
            .I(N__21455));
    InMux I__2556 (
            .O(N__21458),
            .I(N__21452));
    LocalMux I__2555 (
            .O(N__21455),
            .I(N__21447));
    LocalMux I__2554 (
            .O(N__21452),
            .I(N__21447));
    Odrv4 I__2553 (
            .O(N__21447),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2552 (
            .O(N__21444),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    CascadeMux I__2551 (
            .O(N__21441),
            .I(N__21438));
    InMux I__2550 (
            .O(N__21438),
            .I(N__21432));
    InMux I__2549 (
            .O(N__21437),
            .I(N__21429));
    InMux I__2548 (
            .O(N__21436),
            .I(N__21426));
    InMux I__2547 (
            .O(N__21435),
            .I(N__21423));
    LocalMux I__2546 (
            .O(N__21432),
            .I(N__21418));
    LocalMux I__2545 (
            .O(N__21429),
            .I(N__21418));
    LocalMux I__2544 (
            .O(N__21426),
            .I(N__21415));
    LocalMux I__2543 (
            .O(N__21423),
            .I(N__21412));
    Span4Mux_h I__2542 (
            .O(N__21418),
            .I(N__21407));
    Span4Mux_h I__2541 (
            .O(N__21415),
            .I(N__21407));
    Odrv12 I__2540 (
            .O(N__21412),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__2539 (
            .O(N__21407),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__2538 (
            .O(N__21402),
            .I(N__21399));
    LocalMux I__2537 (
            .O(N__21399),
            .I(N__21395));
    InMux I__2536 (
            .O(N__21398),
            .I(N__21392));
    Span4Mux_s3_h I__2535 (
            .O(N__21395),
            .I(N__21387));
    LocalMux I__2534 (
            .O(N__21392),
            .I(N__21387));
    Odrv4 I__2533 (
            .O(N__21387),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2532 (
            .O(N__21384),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2531 (
            .O(N__21381),
            .I(N__21378));
    LocalMux I__2530 (
            .O(N__21378),
            .I(N__21375));
    Odrv12 I__2529 (
            .O(N__21375),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__2528 (
            .O(N__21372),
            .I(N__21367));
    InMux I__2527 (
            .O(N__21371),
            .I(N__21364));
    InMux I__2526 (
            .O(N__21370),
            .I(N__21361));
    InMux I__2525 (
            .O(N__21367),
            .I(N__21357));
    LocalMux I__2524 (
            .O(N__21364),
            .I(N__21354));
    LocalMux I__2523 (
            .O(N__21361),
            .I(N__21351));
    InMux I__2522 (
            .O(N__21360),
            .I(N__21348));
    LocalMux I__2521 (
            .O(N__21357),
            .I(N__21345));
    Span4Mux_s3_h I__2520 (
            .O(N__21354),
            .I(N__21340));
    Span4Mux_s3_h I__2519 (
            .O(N__21351),
            .I(N__21340));
    LocalMux I__2518 (
            .O(N__21348),
            .I(N__21337));
    Odrv4 I__2517 (
            .O(N__21345),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__2516 (
            .O(N__21340),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__2515 (
            .O(N__21337),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__2514 (
            .O(N__21330),
            .I(N__21327));
    InMux I__2513 (
            .O(N__21327),
            .I(N__21323));
    InMux I__2512 (
            .O(N__21326),
            .I(N__21320));
    LocalMux I__2511 (
            .O(N__21323),
            .I(N__21317));
    LocalMux I__2510 (
            .O(N__21320),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    Odrv4 I__2509 (
            .O(N__21317),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2508 (
            .O(N__21312),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2507 (
            .O(N__21309),
            .I(N__21305));
    InMux I__2506 (
            .O(N__21308),
            .I(N__21302));
    LocalMux I__2505 (
            .O(N__21305),
            .I(N__21297));
    LocalMux I__2504 (
            .O(N__21302),
            .I(N__21294));
    InMux I__2503 (
            .O(N__21301),
            .I(N__21291));
    InMux I__2502 (
            .O(N__21300),
            .I(N__21288));
    Span4Mux_h I__2501 (
            .O(N__21297),
            .I(N__21283));
    Span4Mux_h I__2500 (
            .O(N__21294),
            .I(N__21283));
    LocalMux I__2499 (
            .O(N__21291),
            .I(N__21278));
    LocalMux I__2498 (
            .O(N__21288),
            .I(N__21278));
    Odrv4 I__2497 (
            .O(N__21283),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__2496 (
            .O(N__21278),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__2495 (
            .O(N__21273),
            .I(N__21269));
    InMux I__2494 (
            .O(N__21272),
            .I(N__21266));
    LocalMux I__2493 (
            .O(N__21269),
            .I(N__21263));
    LocalMux I__2492 (
            .O(N__21266),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    Odrv4 I__2491 (
            .O(N__21263),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2490 (
            .O(N__21258),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    CascadeMux I__2489 (
            .O(N__21255),
            .I(N__21252));
    InMux I__2488 (
            .O(N__21252),
            .I(N__21248));
    InMux I__2487 (
            .O(N__21251),
            .I(N__21244));
    LocalMux I__2486 (
            .O(N__21248),
            .I(N__21240));
    InMux I__2485 (
            .O(N__21247),
            .I(N__21237));
    LocalMux I__2484 (
            .O(N__21244),
            .I(N__21234));
    InMux I__2483 (
            .O(N__21243),
            .I(N__21231));
    Span4Mux_v I__2482 (
            .O(N__21240),
            .I(N__21228));
    LocalMux I__2481 (
            .O(N__21237),
            .I(N__21225));
    Sp12to4 I__2480 (
            .O(N__21234),
            .I(N__21220));
    LocalMux I__2479 (
            .O(N__21231),
            .I(N__21220));
    Odrv4 I__2478 (
            .O(N__21228),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__2477 (
            .O(N__21225),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv12 I__2476 (
            .O(N__21220),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__2475 (
            .O(N__21213),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    CascadeMux I__2474 (
            .O(N__21210),
            .I(N__21205));
    InMux I__2473 (
            .O(N__21209),
            .I(N__21202));
    InMux I__2472 (
            .O(N__21208),
            .I(N__21199));
    InMux I__2471 (
            .O(N__21205),
            .I(N__21196));
    LocalMux I__2470 (
            .O(N__21202),
            .I(N__21192));
    LocalMux I__2469 (
            .O(N__21199),
            .I(N__21189));
    LocalMux I__2468 (
            .O(N__21196),
            .I(N__21186));
    InMux I__2467 (
            .O(N__21195),
            .I(N__21183));
    Span4Mux_v I__2466 (
            .O(N__21192),
            .I(N__21180));
    Span4Mux_v I__2465 (
            .O(N__21189),
            .I(N__21175));
    Span4Mux_v I__2464 (
            .O(N__21186),
            .I(N__21175));
    LocalMux I__2463 (
            .O(N__21183),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__2462 (
            .O(N__21180),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__2461 (
            .O(N__21175),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__2460 (
            .O(N__21168),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    CascadeMux I__2459 (
            .O(N__21165),
            .I(N__21162));
    InMux I__2458 (
            .O(N__21162),
            .I(N__21157));
    CascadeMux I__2457 (
            .O(N__21161),
            .I(N__21154));
    InMux I__2456 (
            .O(N__21160),
            .I(N__21151));
    LocalMux I__2455 (
            .O(N__21157),
            .I(N__21148));
    InMux I__2454 (
            .O(N__21154),
            .I(N__21145));
    LocalMux I__2453 (
            .O(N__21151),
            .I(N__21142));
    Span4Mux_h I__2452 (
            .O(N__21148),
            .I(N__21136));
    LocalMux I__2451 (
            .O(N__21145),
            .I(N__21136));
    Span4Mux_v I__2450 (
            .O(N__21142),
            .I(N__21133));
    InMux I__2449 (
            .O(N__21141),
            .I(N__21130));
    Span4Mux_v I__2448 (
            .O(N__21136),
            .I(N__21127));
    Odrv4 I__2447 (
            .O(N__21133),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__2446 (
            .O(N__21130),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__2445 (
            .O(N__21127),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__2444 (
            .O(N__21120),
            .I(bfn_3_19_0_));
    InMux I__2443 (
            .O(N__21117),
            .I(N__21114));
    LocalMux I__2442 (
            .O(N__21114),
            .I(N__21111));
    Odrv12 I__2441 (
            .O(N__21111),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__2440 (
            .O(N__21108),
            .I(N__21103));
    InMux I__2439 (
            .O(N__21107),
            .I(N__21098));
    InMux I__2438 (
            .O(N__21106),
            .I(N__21098));
    InMux I__2437 (
            .O(N__21103),
            .I(N__21095));
    LocalMux I__2436 (
            .O(N__21098),
            .I(N__21091));
    LocalMux I__2435 (
            .O(N__21095),
            .I(N__21088));
    CascadeMux I__2434 (
            .O(N__21094),
            .I(N__21085));
    Span4Mux_v I__2433 (
            .O(N__21091),
            .I(N__21082));
    Span4Mux_v I__2432 (
            .O(N__21088),
            .I(N__21079));
    InMux I__2431 (
            .O(N__21085),
            .I(N__21076));
    Odrv4 I__2430 (
            .O(N__21082),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__2429 (
            .O(N__21079),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__2428 (
            .O(N__21076),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__2427 (
            .O(N__21069),
            .I(N__21066));
    LocalMux I__2426 (
            .O(N__21066),
            .I(N__21061));
    InMux I__2425 (
            .O(N__21065),
            .I(N__21056));
    InMux I__2424 (
            .O(N__21064),
            .I(N__21056));
    Span4Mux_v I__2423 (
            .O(N__21061),
            .I(N__21051));
    LocalMux I__2422 (
            .O(N__21056),
            .I(N__21051));
    Span4Mux_v I__2421 (
            .O(N__21051),
            .I(N__21048));
    Odrv4 I__2420 (
            .O(N__21048),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2419 (
            .O(N__21045),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__2418 (
            .O(N__21042),
            .I(N__21039));
    LocalMux I__2417 (
            .O(N__21039),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__2416 (
            .O(N__21036),
            .I(N__21031));
    InMux I__2415 (
            .O(N__21035),
            .I(N__21026));
    InMux I__2414 (
            .O(N__21034),
            .I(N__21026));
    InMux I__2413 (
            .O(N__21031),
            .I(N__21023));
    LocalMux I__2412 (
            .O(N__21026),
            .I(N__21017));
    LocalMux I__2411 (
            .O(N__21023),
            .I(N__21017));
    InMux I__2410 (
            .O(N__21022),
            .I(N__21014));
    Span4Mux_h I__2409 (
            .O(N__21017),
            .I(N__21011));
    LocalMux I__2408 (
            .O(N__21014),
            .I(N__21008));
    Odrv4 I__2407 (
            .O(N__21011),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__2406 (
            .O(N__21008),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__2405 (
            .O(N__21003),
            .I(N__20999));
    InMux I__2404 (
            .O(N__21002),
            .I(N__20996));
    LocalMux I__2403 (
            .O(N__20999),
            .I(N__20989));
    LocalMux I__2402 (
            .O(N__20996),
            .I(N__20989));
    InMux I__2401 (
            .O(N__20995),
            .I(N__20984));
    InMux I__2400 (
            .O(N__20994),
            .I(N__20984));
    Span4Mux_v I__2399 (
            .O(N__20989),
            .I(N__20979));
    LocalMux I__2398 (
            .O(N__20984),
            .I(N__20979));
    Span4Mux_v I__2397 (
            .O(N__20979),
            .I(N__20976));
    Odrv4 I__2396 (
            .O(N__20976),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2395 (
            .O(N__20973),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2394 (
            .O(N__20970),
            .I(N__20967));
    LocalMux I__2393 (
            .O(N__20967),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__2392 (
            .O(N__20964),
            .I(N__20961));
    InMux I__2391 (
            .O(N__20961),
            .I(N__20958));
    LocalMux I__2390 (
            .O(N__20958),
            .I(N__20953));
    InMux I__2389 (
            .O(N__20957),
            .I(N__20948));
    InMux I__2388 (
            .O(N__20956),
            .I(N__20948));
    Span4Mux_h I__2387 (
            .O(N__20953),
            .I(N__20943));
    LocalMux I__2386 (
            .O(N__20948),
            .I(N__20943));
    Span4Mux_v I__2385 (
            .O(N__20943),
            .I(N__20939));
    InMux I__2384 (
            .O(N__20942),
            .I(N__20936));
    Odrv4 I__2383 (
            .O(N__20939),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__2382 (
            .O(N__20936),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__2381 (
            .O(N__20931),
            .I(N__20928));
    LocalMux I__2380 (
            .O(N__20928),
            .I(N__20923));
    InMux I__2379 (
            .O(N__20927),
            .I(N__20920));
    CascadeMux I__2378 (
            .O(N__20926),
            .I(N__20917));
    Span4Mux_v I__2377 (
            .O(N__20923),
            .I(N__20914));
    LocalMux I__2376 (
            .O(N__20920),
            .I(N__20911));
    InMux I__2375 (
            .O(N__20917),
            .I(N__20908));
    Span4Mux_v I__2374 (
            .O(N__20914),
            .I(N__20905));
    Span4Mux_v I__2373 (
            .O(N__20911),
            .I(N__20900));
    LocalMux I__2372 (
            .O(N__20908),
            .I(N__20900));
    Odrv4 I__2371 (
            .O(N__20905),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__2370 (
            .O(N__20900),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2369 (
            .O(N__20895),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2368 (
            .O(N__20892),
            .I(N__20889));
    LocalMux I__2367 (
            .O(N__20889),
            .I(N__20886));
    Odrv4 I__2366 (
            .O(N__20886),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__2365 (
            .O(N__20883),
            .I(N__20879));
    CascadeMux I__2364 (
            .O(N__20882),
            .I(N__20875));
    InMux I__2363 (
            .O(N__20879),
            .I(N__20872));
    InMux I__2362 (
            .O(N__20878),
            .I(N__20869));
    InMux I__2361 (
            .O(N__20875),
            .I(N__20866));
    LocalMux I__2360 (
            .O(N__20872),
            .I(N__20863));
    LocalMux I__2359 (
            .O(N__20869),
            .I(N__20857));
    LocalMux I__2358 (
            .O(N__20866),
            .I(N__20857));
    Span4Mux_v I__2357 (
            .O(N__20863),
            .I(N__20854));
    InMux I__2356 (
            .O(N__20862),
            .I(N__20851));
    Odrv12 I__2355 (
            .O(N__20857),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__2354 (
            .O(N__20854),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__2353 (
            .O(N__20851),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__2352 (
            .O(N__20844),
            .I(N__20841));
    LocalMux I__2351 (
            .O(N__20841),
            .I(N__20837));
    InMux I__2350 (
            .O(N__20840),
            .I(N__20834));
    Span4Mux_s3_h I__2349 (
            .O(N__20837),
            .I(N__20830));
    LocalMux I__2348 (
            .O(N__20834),
            .I(N__20827));
    InMux I__2347 (
            .O(N__20833),
            .I(N__20824));
    Span4Mux_v I__2346 (
            .O(N__20830),
            .I(N__20821));
    Span4Mux_v I__2345 (
            .O(N__20827),
            .I(N__20816));
    LocalMux I__2344 (
            .O(N__20824),
            .I(N__20816));
    Odrv4 I__2343 (
            .O(N__20821),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2342 (
            .O(N__20816),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2341 (
            .O(N__20811),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__2340 (
            .O(N__20808),
            .I(N__20805));
    LocalMux I__2339 (
            .O(N__20805),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__2338 (
            .O(N__20802),
            .I(N__20799));
    InMux I__2337 (
            .O(N__20799),
            .I(N__20796));
    LocalMux I__2336 (
            .O(N__20796),
            .I(N__20792));
    InMux I__2335 (
            .O(N__20795),
            .I(N__20787));
    Span4Mux_h I__2334 (
            .O(N__20792),
            .I(N__20784));
    InMux I__2333 (
            .O(N__20791),
            .I(N__20779));
    InMux I__2332 (
            .O(N__20790),
            .I(N__20779));
    LocalMux I__2331 (
            .O(N__20787),
            .I(N__20776));
    Odrv4 I__2330 (
            .O(N__20784),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__2329 (
            .O(N__20779),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv12 I__2328 (
            .O(N__20776),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    CascadeMux I__2327 (
            .O(N__20769),
            .I(N__20766));
    InMux I__2326 (
            .O(N__20766),
            .I(N__20761));
    InMux I__2325 (
            .O(N__20765),
            .I(N__20758));
    InMux I__2324 (
            .O(N__20764),
            .I(N__20755));
    LocalMux I__2323 (
            .O(N__20761),
            .I(N__20752));
    LocalMux I__2322 (
            .O(N__20758),
            .I(N__20749));
    LocalMux I__2321 (
            .O(N__20755),
            .I(N__20746));
    Span12Mux_s3_h I__2320 (
            .O(N__20752),
            .I(N__20743));
    Span4Mux_v I__2319 (
            .O(N__20749),
            .I(N__20738));
    Span4Mux_s3_h I__2318 (
            .O(N__20746),
            .I(N__20738));
    Odrv12 I__2317 (
            .O(N__20743),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2316 (
            .O(N__20738),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2315 (
            .O(N__20733),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    CascadeMux I__2314 (
            .O(N__20730),
            .I(N__20724));
    InMux I__2313 (
            .O(N__20729),
            .I(N__20719));
    InMux I__2312 (
            .O(N__20728),
            .I(N__20719));
    InMux I__2311 (
            .O(N__20727),
            .I(N__20716));
    InMux I__2310 (
            .O(N__20724),
            .I(N__20713));
    LocalMux I__2309 (
            .O(N__20719),
            .I(N__20710));
    LocalMux I__2308 (
            .O(N__20716),
            .I(N__20707));
    LocalMux I__2307 (
            .O(N__20713),
            .I(N__20704));
    Span4Mux_v I__2306 (
            .O(N__20710),
            .I(N__20701));
    Span4Mux_s3_h I__2305 (
            .O(N__20707),
            .I(N__20698));
    Odrv12 I__2304 (
            .O(N__20704),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__2303 (
            .O(N__20701),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__2302 (
            .O(N__20698),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__2301 (
            .O(N__20691),
            .I(N__20688));
    LocalMux I__2300 (
            .O(N__20688),
            .I(N__20684));
    InMux I__2299 (
            .O(N__20687),
            .I(N__20680));
    Span4Mux_h I__2298 (
            .O(N__20684),
            .I(N__20677));
    InMux I__2297 (
            .O(N__20683),
            .I(N__20674));
    LocalMux I__2296 (
            .O(N__20680),
            .I(N__20671));
    Span4Mux_v I__2295 (
            .O(N__20677),
            .I(N__20668));
    LocalMux I__2294 (
            .O(N__20674),
            .I(N__20663));
    Span4Mux_v I__2293 (
            .O(N__20671),
            .I(N__20663));
    Odrv4 I__2292 (
            .O(N__20668),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2291 (
            .O(N__20663),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2290 (
            .O(N__20658),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    CascadeMux I__2289 (
            .O(N__20655),
            .I(N__20651));
    CascadeMux I__2288 (
            .O(N__20654),
            .I(N__20648));
    InMux I__2287 (
            .O(N__20651),
            .I(N__20643));
    InMux I__2286 (
            .O(N__20648),
            .I(N__20640));
    InMux I__2285 (
            .O(N__20647),
            .I(N__20635));
    InMux I__2284 (
            .O(N__20646),
            .I(N__20635));
    LocalMux I__2283 (
            .O(N__20643),
            .I(N__20632));
    LocalMux I__2282 (
            .O(N__20640),
            .I(N__20629));
    LocalMux I__2281 (
            .O(N__20635),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__2280 (
            .O(N__20632),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__2279 (
            .O(N__20629),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    CascadeMux I__2278 (
            .O(N__20622),
            .I(N__20619));
    InMux I__2277 (
            .O(N__20619),
            .I(N__20616));
    LocalMux I__2276 (
            .O(N__20616),
            .I(N__20612));
    InMux I__2275 (
            .O(N__20615),
            .I(N__20609));
    Span4Mux_s3_h I__2274 (
            .O(N__20612),
            .I(N__20605));
    LocalMux I__2273 (
            .O(N__20609),
            .I(N__20602));
    InMux I__2272 (
            .O(N__20608),
            .I(N__20599));
    Span4Mux_v I__2271 (
            .O(N__20605),
            .I(N__20596));
    Span4Mux_v I__2270 (
            .O(N__20602),
            .I(N__20591));
    LocalMux I__2269 (
            .O(N__20599),
            .I(N__20591));
    Odrv4 I__2268 (
            .O(N__20596),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__2267 (
            .O(N__20591),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2266 (
            .O(N__20586),
            .I(bfn_3_18_0_));
    InMux I__2265 (
            .O(N__20583),
            .I(N__20580));
    LocalMux I__2264 (
            .O(N__20580),
            .I(N__20577));
    Span4Mux_v I__2263 (
            .O(N__20577),
            .I(N__20574));
    Span4Mux_v I__2262 (
            .O(N__20574),
            .I(N__20571));
    Odrv4 I__2261 (
            .O(N__20571),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2260 (
            .O(N__20568),
            .I(N__20562));
    InMux I__2259 (
            .O(N__20567),
            .I(N__20548));
    InMux I__2258 (
            .O(N__20566),
            .I(N__20545));
    InMux I__2257 (
            .O(N__20565),
            .I(N__20542));
    LocalMux I__2256 (
            .O(N__20562),
            .I(N__20539));
    InMux I__2255 (
            .O(N__20561),
            .I(N__20536));
    CascadeMux I__2254 (
            .O(N__20560),
            .I(N__20533));
    CascadeMux I__2253 (
            .O(N__20559),
            .I(N__20530));
    CascadeMux I__2252 (
            .O(N__20558),
            .I(N__20527));
    InMux I__2251 (
            .O(N__20557),
            .I(N__20508));
    InMux I__2250 (
            .O(N__20556),
            .I(N__20505));
    InMux I__2249 (
            .O(N__20555),
            .I(N__20494));
    InMux I__2248 (
            .O(N__20554),
            .I(N__20494));
    InMux I__2247 (
            .O(N__20553),
            .I(N__20494));
    InMux I__2246 (
            .O(N__20552),
            .I(N__20494));
    InMux I__2245 (
            .O(N__20551),
            .I(N__20494));
    LocalMux I__2244 (
            .O(N__20548),
            .I(N__20483));
    LocalMux I__2243 (
            .O(N__20545),
            .I(N__20483));
    LocalMux I__2242 (
            .O(N__20542),
            .I(N__20483));
    Span4Mux_h I__2241 (
            .O(N__20539),
            .I(N__20483));
    LocalMux I__2240 (
            .O(N__20536),
            .I(N__20483));
    InMux I__2239 (
            .O(N__20533),
            .I(N__20470));
    InMux I__2238 (
            .O(N__20530),
            .I(N__20470));
    InMux I__2237 (
            .O(N__20527),
            .I(N__20470));
    InMux I__2236 (
            .O(N__20526),
            .I(N__20470));
    InMux I__2235 (
            .O(N__20525),
            .I(N__20470));
    InMux I__2234 (
            .O(N__20524),
            .I(N__20470));
    InMux I__2233 (
            .O(N__20523),
            .I(N__20467));
    InMux I__2232 (
            .O(N__20522),
            .I(N__20452));
    InMux I__2231 (
            .O(N__20521),
            .I(N__20452));
    InMux I__2230 (
            .O(N__20520),
            .I(N__20452));
    InMux I__2229 (
            .O(N__20519),
            .I(N__20452));
    InMux I__2228 (
            .O(N__20518),
            .I(N__20452));
    InMux I__2227 (
            .O(N__20517),
            .I(N__20452));
    InMux I__2226 (
            .O(N__20516),
            .I(N__20452));
    InMux I__2225 (
            .O(N__20515),
            .I(N__20441));
    InMux I__2224 (
            .O(N__20514),
            .I(N__20441));
    InMux I__2223 (
            .O(N__20513),
            .I(N__20441));
    InMux I__2222 (
            .O(N__20512),
            .I(N__20441));
    InMux I__2221 (
            .O(N__20511),
            .I(N__20441));
    LocalMux I__2220 (
            .O(N__20508),
            .I(N__20434));
    LocalMux I__2219 (
            .O(N__20505),
            .I(N__20434));
    LocalMux I__2218 (
            .O(N__20494),
            .I(N__20434));
    Span4Mux_v I__2217 (
            .O(N__20483),
            .I(N__20431));
    LocalMux I__2216 (
            .O(N__20470),
            .I(N__20422));
    LocalMux I__2215 (
            .O(N__20467),
            .I(N__20422));
    LocalMux I__2214 (
            .O(N__20452),
            .I(N__20422));
    LocalMux I__2213 (
            .O(N__20441),
            .I(N__20422));
    Odrv4 I__2212 (
            .O(N__20434),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2211 (
            .O(N__20431),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv12 I__2210 (
            .O(N__20422),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    CascadeMux I__2209 (
            .O(N__20415),
            .I(N__20412));
    InMux I__2208 (
            .O(N__20412),
            .I(N__20409));
    LocalMux I__2207 (
            .O(N__20409),
            .I(N__20406));
    Span4Mux_h I__2206 (
            .O(N__20406),
            .I(N__20403));
    Odrv4 I__2205 (
            .O(N__20403),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    CascadeMux I__2204 (
            .O(N__20400),
            .I(N__20391));
    CascadeMux I__2203 (
            .O(N__20399),
            .I(N__20388));
    InMux I__2202 (
            .O(N__20398),
            .I(N__20382));
    InMux I__2201 (
            .O(N__20397),
            .I(N__20379));
    InMux I__2200 (
            .O(N__20396),
            .I(N__20357));
    InMux I__2199 (
            .O(N__20395),
            .I(N__20357));
    InMux I__2198 (
            .O(N__20394),
            .I(N__20357));
    InMux I__2197 (
            .O(N__20391),
            .I(N__20357));
    InMux I__2196 (
            .O(N__20388),
            .I(N__20357));
    InMux I__2195 (
            .O(N__20387),
            .I(N__20347));
    InMux I__2194 (
            .O(N__20386),
            .I(N__20344));
    InMux I__2193 (
            .O(N__20385),
            .I(N__20341));
    LocalMux I__2192 (
            .O(N__20382),
            .I(N__20336));
    LocalMux I__2191 (
            .O(N__20379),
            .I(N__20336));
    InMux I__2190 (
            .O(N__20378),
            .I(N__20333));
    InMux I__2189 (
            .O(N__20377),
            .I(N__20326));
    InMux I__2188 (
            .O(N__20376),
            .I(N__20326));
    InMux I__2187 (
            .O(N__20375),
            .I(N__20326));
    InMux I__2186 (
            .O(N__20374),
            .I(N__20317));
    InMux I__2185 (
            .O(N__20373),
            .I(N__20317));
    InMux I__2184 (
            .O(N__20372),
            .I(N__20317));
    InMux I__2183 (
            .O(N__20371),
            .I(N__20317));
    CascadeMux I__2182 (
            .O(N__20370),
            .I(N__20311));
    CascadeMux I__2181 (
            .O(N__20369),
            .I(N__20308));
    CascadeMux I__2180 (
            .O(N__20368),
            .I(N__20305));
    LocalMux I__2179 (
            .O(N__20357),
            .I(N__20302));
    InMux I__2178 (
            .O(N__20356),
            .I(N__20287));
    InMux I__2177 (
            .O(N__20355),
            .I(N__20287));
    InMux I__2176 (
            .O(N__20354),
            .I(N__20287));
    InMux I__2175 (
            .O(N__20353),
            .I(N__20287));
    InMux I__2174 (
            .O(N__20352),
            .I(N__20287));
    InMux I__2173 (
            .O(N__20351),
            .I(N__20287));
    InMux I__2172 (
            .O(N__20350),
            .I(N__20287));
    LocalMux I__2171 (
            .O(N__20347),
            .I(N__20282));
    LocalMux I__2170 (
            .O(N__20344),
            .I(N__20282));
    LocalMux I__2169 (
            .O(N__20341),
            .I(N__20277));
    Span4Mux_v I__2168 (
            .O(N__20336),
            .I(N__20277));
    LocalMux I__2167 (
            .O(N__20333),
            .I(N__20274));
    LocalMux I__2166 (
            .O(N__20326),
            .I(N__20269));
    LocalMux I__2165 (
            .O(N__20317),
            .I(N__20269));
    InMux I__2164 (
            .O(N__20316),
            .I(N__20266));
    InMux I__2163 (
            .O(N__20315),
            .I(N__20255));
    InMux I__2162 (
            .O(N__20314),
            .I(N__20255));
    InMux I__2161 (
            .O(N__20311),
            .I(N__20255));
    InMux I__2160 (
            .O(N__20308),
            .I(N__20255));
    InMux I__2159 (
            .O(N__20305),
            .I(N__20255));
    Span4Mux_h I__2158 (
            .O(N__20302),
            .I(N__20250));
    LocalMux I__2157 (
            .O(N__20287),
            .I(N__20250));
    Span4Mux_v I__2156 (
            .O(N__20282),
            .I(N__20245));
    Span4Mux_v I__2155 (
            .O(N__20277),
            .I(N__20245));
    Span4Mux_v I__2154 (
            .O(N__20274),
            .I(N__20240));
    Span4Mux_v I__2153 (
            .O(N__20269),
            .I(N__20240));
    LocalMux I__2152 (
            .O(N__20266),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    LocalMux I__2151 (
            .O(N__20255),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2150 (
            .O(N__20250),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2149 (
            .O(N__20245),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2148 (
            .O(N__20240),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    InMux I__2147 (
            .O(N__20229),
            .I(N__20225));
    InMux I__2146 (
            .O(N__20228),
            .I(N__20222));
    LocalMux I__2145 (
            .O(N__20225),
            .I(N__20219));
    LocalMux I__2144 (
            .O(N__20222),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    Odrv4 I__2143 (
            .O(N__20219),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__2142 (
            .O(N__20214),
            .I(N__20210));
    InMux I__2141 (
            .O(N__20213),
            .I(N__20206));
    InMux I__2140 (
            .O(N__20210),
            .I(N__20203));
    CascadeMux I__2139 (
            .O(N__20209),
            .I(N__20200));
    LocalMux I__2138 (
            .O(N__20206),
            .I(N__20195));
    LocalMux I__2137 (
            .O(N__20203),
            .I(N__20195));
    InMux I__2136 (
            .O(N__20200),
            .I(N__20191));
    Span4Mux_v I__2135 (
            .O(N__20195),
            .I(N__20188));
    InMux I__2134 (
            .O(N__20194),
            .I(N__20184));
    LocalMux I__2133 (
            .O(N__20191),
            .I(N__20181));
    Span4Mux_s3_h I__2132 (
            .O(N__20188),
            .I(N__20178));
    InMux I__2131 (
            .O(N__20187),
            .I(N__20175));
    LocalMux I__2130 (
            .O(N__20184),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__2129 (
            .O(N__20181),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__2128 (
            .O(N__20178),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__2127 (
            .O(N__20175),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__2126 (
            .O(N__20166),
            .I(N__20162));
    InMux I__2125 (
            .O(N__20165),
            .I(N__20159));
    InMux I__2124 (
            .O(N__20162),
            .I(N__20156));
    LocalMux I__2123 (
            .O(N__20159),
            .I(N__20152));
    LocalMux I__2122 (
            .O(N__20156),
            .I(N__20149));
    InMux I__2121 (
            .O(N__20155),
            .I(N__20146));
    Span4Mux_v I__2120 (
            .O(N__20152),
            .I(N__20143));
    Span4Mux_v I__2119 (
            .O(N__20149),
            .I(N__20140));
    LocalMux I__2118 (
            .O(N__20146),
            .I(N__20137));
    Odrv4 I__2117 (
            .O(N__20143),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__2116 (
            .O(N__20140),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__2115 (
            .O(N__20137),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__2114 (
            .O(N__20130),
            .I(N__20127));
    LocalMux I__2113 (
            .O(N__20127),
            .I(N__20124));
    Span4Mux_h I__2112 (
            .O(N__20124),
            .I(N__20121));
    Span4Mux_v I__2111 (
            .O(N__20121),
            .I(N__20118));
    Odrv4 I__2110 (
            .O(N__20118),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2109 (
            .O(N__20115),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2108 (
            .O(N__20112),
            .I(N__20109));
    LocalMux I__2107 (
            .O(N__20109),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    InMux I__2106 (
            .O(N__20106),
            .I(N__20102));
    InMux I__2105 (
            .O(N__20105),
            .I(N__20098));
    LocalMux I__2104 (
            .O(N__20102),
            .I(N__20095));
    InMux I__2103 (
            .O(N__20101),
            .I(N__20092));
    LocalMux I__2102 (
            .O(N__20098),
            .I(N__20089));
    Odrv4 I__2101 (
            .O(N__20095),
            .I(pwm_duty_input_4));
    LocalMux I__2100 (
            .O(N__20092),
            .I(pwm_duty_input_4));
    Odrv4 I__2099 (
            .O(N__20089),
            .I(pwm_duty_input_4));
    CascadeMux I__2098 (
            .O(N__20082),
            .I(N__20079));
    InMux I__2097 (
            .O(N__20079),
            .I(N__20075));
    InMux I__2096 (
            .O(N__20078),
            .I(N__20071));
    LocalMux I__2095 (
            .O(N__20075),
            .I(N__20068));
    InMux I__2094 (
            .O(N__20074),
            .I(N__20065));
    LocalMux I__2093 (
            .O(N__20071),
            .I(N__20062));
    Odrv4 I__2092 (
            .O(N__20068),
            .I(pwm_duty_input_3));
    LocalMux I__2091 (
            .O(N__20065),
            .I(pwm_duty_input_3));
    Odrv4 I__2090 (
            .O(N__20062),
            .I(pwm_duty_input_3));
    InMux I__2089 (
            .O(N__20055),
            .I(N__20051));
    InMux I__2088 (
            .O(N__20054),
            .I(N__20048));
    LocalMux I__2087 (
            .O(N__20051),
            .I(N__20044));
    LocalMux I__2086 (
            .O(N__20048),
            .I(N__20041));
    InMux I__2085 (
            .O(N__20047),
            .I(N__20038));
    Span4Mux_v I__2084 (
            .O(N__20044),
            .I(N__20035));
    Odrv4 I__2083 (
            .O(N__20041),
            .I(pwm_duty_input_5));
    LocalMux I__2082 (
            .O(N__20038),
            .I(pwm_duty_input_5));
    Odrv4 I__2081 (
            .O(N__20035),
            .I(pwm_duty_input_5));
    InMux I__2080 (
            .O(N__20028),
            .I(N__20025));
    LocalMux I__2079 (
            .O(N__20025),
            .I(N__20022));
    Odrv4 I__2078 (
            .O(N__20022),
            .I(rgb_drv_RNOZ0));
    InMux I__2077 (
            .O(N__20019),
            .I(N__20016));
    LocalMux I__2076 (
            .O(N__20016),
            .I(N__20013));
    Odrv4 I__2075 (
            .O(N__20013),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    CascadeMux I__2074 (
            .O(N__20010),
            .I(N__20007));
    InMux I__2073 (
            .O(N__20007),
            .I(N__20004));
    LocalMux I__2072 (
            .O(N__20004),
            .I(N__20001));
    Span4Mux_h I__2071 (
            .O(N__20001),
            .I(N__19998));
    Odrv4 I__2070 (
            .O(N__19998),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    CascadeMux I__2069 (
            .O(N__19995),
            .I(N__19992));
    InMux I__2068 (
            .O(N__19992),
            .I(N__19989));
    LocalMux I__2067 (
            .O(N__19989),
            .I(N__19986));
    Span4Mux_h I__2066 (
            .O(N__19986),
            .I(N__19983));
    Odrv4 I__2065 (
            .O(N__19983),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    CascadeMux I__2064 (
            .O(N__19980),
            .I(N__19977));
    InMux I__2063 (
            .O(N__19977),
            .I(N__19974));
    LocalMux I__2062 (
            .O(N__19974),
            .I(N__19971));
    Span4Mux_h I__2061 (
            .O(N__19971),
            .I(N__19968));
    Odrv4 I__2060 (
            .O(N__19968),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    CascadeMux I__2059 (
            .O(N__19965),
            .I(N__19957));
    InMux I__2058 (
            .O(N__19964),
            .I(N__19948));
    InMux I__2057 (
            .O(N__19963),
            .I(N__19948));
    InMux I__2056 (
            .O(N__19962),
            .I(N__19948));
    InMux I__2055 (
            .O(N__19961),
            .I(N__19948));
    InMux I__2054 (
            .O(N__19960),
            .I(N__19940));
    InMux I__2053 (
            .O(N__19957),
            .I(N__19940));
    LocalMux I__2052 (
            .O(N__19948),
            .I(N__19937));
    InMux I__2051 (
            .O(N__19947),
            .I(N__19934));
    InMux I__2050 (
            .O(N__19946),
            .I(N__19931));
    InMux I__2049 (
            .O(N__19945),
            .I(N__19928));
    LocalMux I__2048 (
            .O(N__19940),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    Odrv4 I__2047 (
            .O(N__19937),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    LocalMux I__2046 (
            .O(N__19934),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    LocalMux I__2045 (
            .O(N__19931),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    LocalMux I__2044 (
            .O(N__19928),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    CascadeMux I__2043 (
            .O(N__19917),
            .I(N__19914));
    InMux I__2042 (
            .O(N__19914),
            .I(N__19908));
    InMux I__2041 (
            .O(N__19913),
            .I(N__19908));
    LocalMux I__2040 (
            .O(N__19908),
            .I(N__19904));
    InMux I__2039 (
            .O(N__19907),
            .I(N__19901));
    Odrv12 I__2038 (
            .O(N__19904),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__2037 (
            .O(N__19901),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__2036 (
            .O(N__19896),
            .I(N__19893));
    LocalMux I__2035 (
            .O(N__19893),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    CascadeMux I__2034 (
            .O(N__19890),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ));
    InMux I__2033 (
            .O(N__19887),
            .I(N__19883));
    InMux I__2032 (
            .O(N__19886),
            .I(N__19880));
    LocalMux I__2031 (
            .O(N__19883),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__2030 (
            .O(N__19880),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__2029 (
            .O(N__19875),
            .I(N__19872));
    LocalMux I__2028 (
            .O(N__19872),
            .I(N__19868));
    InMux I__2027 (
            .O(N__19871),
            .I(N__19865));
    Span4Mux_v I__2026 (
            .O(N__19868),
            .I(N__19862));
    LocalMux I__2025 (
            .O(N__19865),
            .I(pwm_duty_input_0));
    Odrv4 I__2024 (
            .O(N__19862),
            .I(pwm_duty_input_0));
    InMux I__2023 (
            .O(N__19857),
            .I(N__19853));
    InMux I__2022 (
            .O(N__19856),
            .I(N__19850));
    LocalMux I__2021 (
            .O(N__19853),
            .I(N__19847));
    LocalMux I__2020 (
            .O(N__19850),
            .I(pwm_duty_input_1));
    Odrv4 I__2019 (
            .O(N__19847),
            .I(pwm_duty_input_1));
    InMux I__2018 (
            .O(N__19842),
            .I(N__19839));
    LocalMux I__2017 (
            .O(N__19839),
            .I(N__19835));
    InMux I__2016 (
            .O(N__19838),
            .I(N__19832));
    Span4Mux_s1_h I__2015 (
            .O(N__19835),
            .I(N__19829));
    LocalMux I__2014 (
            .O(N__19832),
            .I(pwm_duty_input_2));
    Odrv4 I__2013 (
            .O(N__19829),
            .I(pwm_duty_input_2));
    InMux I__2012 (
            .O(N__19824),
            .I(N__19819));
    InMux I__2011 (
            .O(N__19823),
            .I(N__19814));
    InMux I__2010 (
            .O(N__19822),
            .I(N__19814));
    LocalMux I__2009 (
            .O(N__19819),
            .I(N__19811));
    LocalMux I__2008 (
            .O(N__19814),
            .I(pwm_duty_input_7));
    Odrv4 I__2007 (
            .O(N__19811),
            .I(pwm_duty_input_7));
    InMux I__2006 (
            .O(N__19806),
            .I(N__19803));
    LocalMux I__2005 (
            .O(N__19803),
            .I(N__19798));
    InMux I__2004 (
            .O(N__19802),
            .I(N__19793));
    InMux I__2003 (
            .O(N__19801),
            .I(N__19793));
    Span4Mux_v I__2002 (
            .O(N__19798),
            .I(N__19790));
    LocalMux I__2001 (
            .O(N__19793),
            .I(pwm_duty_input_8));
    Odrv4 I__2000 (
            .O(N__19790),
            .I(pwm_duty_input_8));
    InMux I__1999 (
            .O(N__19785),
            .I(N__19781));
    CascadeMux I__1998 (
            .O(N__19784),
            .I(N__19777));
    LocalMux I__1997 (
            .O(N__19781),
            .I(N__19774));
    InMux I__1996 (
            .O(N__19780),
            .I(N__19769));
    InMux I__1995 (
            .O(N__19777),
            .I(N__19769));
    Span4Mux_s1_h I__1994 (
            .O(N__19774),
            .I(N__19766));
    LocalMux I__1993 (
            .O(N__19769),
            .I(pwm_duty_input_6));
    Odrv4 I__1992 (
            .O(N__19766),
            .I(pwm_duty_input_6));
    CascadeMux I__1991 (
            .O(N__19761),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__1990 (
            .O(N__19758),
            .I(N__19755));
    LocalMux I__1989 (
            .O(N__19755),
            .I(N__19750));
    InMux I__1988 (
            .O(N__19754),
            .I(N__19745));
    InMux I__1987 (
            .O(N__19753),
            .I(N__19745));
    Span4Mux_s1_h I__1986 (
            .O(N__19750),
            .I(N__19742));
    LocalMux I__1985 (
            .O(N__19745),
            .I(pwm_duty_input_9));
    Odrv4 I__1984 (
            .O(N__19742),
            .I(pwm_duty_input_9));
    InMux I__1983 (
            .O(N__19737),
            .I(N__19734));
    LocalMux I__1982 (
            .O(N__19734),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    CascadeMux I__1981 (
            .O(N__19731),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ));
    CascadeMux I__1980 (
            .O(N__19728),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__1979 (
            .O(N__19725),
            .I(N__19722));
    LocalMux I__1978 (
            .O(N__19722),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__1977 (
            .O(N__19719),
            .I(N__19716));
    LocalMux I__1976 (
            .O(N__19716),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    CascadeMux I__1975 (
            .O(N__19713),
            .I(N__19710));
    InMux I__1974 (
            .O(N__19710),
            .I(N__19707));
    LocalMux I__1973 (
            .O(N__19707),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    CascadeMux I__1972 (
            .O(N__19704),
            .I(N__19696));
    CascadeMux I__1971 (
            .O(N__19703),
            .I(N__19693));
    CascadeMux I__1970 (
            .O(N__19702),
            .I(N__19690));
    CascadeMux I__1969 (
            .O(N__19701),
            .I(N__19687));
    InMux I__1968 (
            .O(N__19700),
            .I(N__19678));
    InMux I__1967 (
            .O(N__19699),
            .I(N__19678));
    InMux I__1966 (
            .O(N__19696),
            .I(N__19678));
    InMux I__1965 (
            .O(N__19693),
            .I(N__19678));
    InMux I__1964 (
            .O(N__19690),
            .I(N__19674));
    InMux I__1963 (
            .O(N__19687),
            .I(N__19671));
    LocalMux I__1962 (
            .O(N__19678),
            .I(N__19668));
    InMux I__1961 (
            .O(N__19677),
            .I(N__19665));
    LocalMux I__1960 (
            .O(N__19674),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    LocalMux I__1959 (
            .O(N__19671),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    Odrv4 I__1958 (
            .O(N__19668),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    LocalMux I__1957 (
            .O(N__19665),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    CascadeMux I__1956 (
            .O(N__19656),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ));
    InMux I__1955 (
            .O(N__19653),
            .I(N__19650));
    LocalMux I__1954 (
            .O(N__19650),
            .I(N__19647));
    Odrv4 I__1953 (
            .O(N__19647),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__1952 (
            .O(N__19644),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ));
    InMux I__1951 (
            .O(N__19641),
            .I(N__19632));
    InMux I__1950 (
            .O(N__19640),
            .I(N__19632));
    InMux I__1949 (
            .O(N__19639),
            .I(N__19632));
    LocalMux I__1948 (
            .O(N__19632),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    CascadeMux I__1947 (
            .O(N__19629),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    CascadeMux I__1946 (
            .O(N__19626),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ));
    InMux I__1945 (
            .O(N__19623),
            .I(N__19620));
    LocalMux I__1944 (
            .O(N__19620),
            .I(\current_shift_inst.PI_CTRL.N_44 ));
    InMux I__1943 (
            .O(N__19617),
            .I(N__19614));
    LocalMux I__1942 (
            .O(N__19614),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    CascadeMux I__1941 (
            .O(N__19611),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_ ));
    InMux I__1940 (
            .O(N__19608),
            .I(N__19605));
    LocalMux I__1939 (
            .O(N__19605),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ));
    InMux I__1938 (
            .O(N__19602),
            .I(N__19599));
    LocalMux I__1937 (
            .O(N__19599),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    CascadeMux I__1936 (
            .O(N__19596),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__1935 (
            .O(N__19593),
            .I(N__19590));
    LocalMux I__1934 (
            .O(N__19590),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    CascadeMux I__1933 (
            .O(N__19587),
            .I(N__19584));
    InMux I__1932 (
            .O(N__19584),
            .I(N__19581));
    LocalMux I__1931 (
            .O(N__19581),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__1930 (
            .O(N__19578),
            .I(N__19575));
    LocalMux I__1929 (
            .O(N__19575),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    CascadeMux I__1928 (
            .O(N__19572),
            .I(N__19569));
    InMux I__1927 (
            .O(N__19569),
            .I(N__19566));
    LocalMux I__1926 (
            .O(N__19566),
            .I(N__19563));
    Span4Mux_v I__1925 (
            .O(N__19563),
            .I(N__19560));
    Odrv4 I__1924 (
            .O(N__19560),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    CascadeMux I__1923 (
            .O(N__19557),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ));
    CascadeMux I__1922 (
            .O(N__19554),
            .I(\current_shift_inst.PI_CTRL.N_77_cascade_ ));
    InMux I__1921 (
            .O(N__19551),
            .I(N__19548));
    LocalMux I__1920 (
            .O(N__19548),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    InMux I__1919 (
            .O(N__19545),
            .I(N__19542));
    LocalMux I__1918 (
            .O(N__19542),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ));
    InMux I__1917 (
            .O(N__19539),
            .I(N__19536));
    LocalMux I__1916 (
            .O(N__19536),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    CascadeMux I__1915 (
            .O(N__19533),
            .I(N__19530));
    InMux I__1914 (
            .O(N__19530),
            .I(N__19527));
    LocalMux I__1913 (
            .O(N__19527),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__1912 (
            .O(N__19524),
            .I(N__19521));
    LocalMux I__1911 (
            .O(N__19521),
            .I(N__19518));
    Odrv4 I__1910 (
            .O(N__19518),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    CascadeMux I__1909 (
            .O(N__19515),
            .I(N__19512));
    InMux I__1908 (
            .O(N__19512),
            .I(N__19509));
    LocalMux I__1907 (
            .O(N__19509),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    CascadeMux I__1906 (
            .O(N__19506),
            .I(N__19503));
    InMux I__1905 (
            .O(N__19503),
            .I(N__19500));
    LocalMux I__1904 (
            .O(N__19500),
            .I(N__19497));
    Odrv4 I__1903 (
            .O(N__19497),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    CascadeMux I__1902 (
            .O(N__19494),
            .I(N__19491));
    InMux I__1901 (
            .O(N__19491),
            .I(N__19488));
    LocalMux I__1900 (
            .O(N__19488),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    CascadeMux I__1899 (
            .O(N__19485),
            .I(N__19482));
    InMux I__1898 (
            .O(N__19482),
            .I(N__19479));
    LocalMux I__1897 (
            .O(N__19479),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    CascadeMux I__1896 (
            .O(N__19476),
            .I(N__19473));
    InMux I__1895 (
            .O(N__19473),
            .I(N__19470));
    LocalMux I__1894 (
            .O(N__19470),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__1893 (
            .O(N__19467),
            .I(N__19464));
    LocalMux I__1892 (
            .O(N__19464),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__1891 (
            .O(N__19461),
            .I(N__19458));
    LocalMux I__1890 (
            .O(N__19458),
            .I(N_38_i_i));
    CascadeMux I__1889 (
            .O(N__19455),
            .I(N__19451));
    CascadeMux I__1888 (
            .O(N__19454),
            .I(N__19448));
    InMux I__1887 (
            .O(N__19451),
            .I(N__19445));
    InMux I__1886 (
            .O(N__19448),
            .I(N__19442));
    LocalMux I__1885 (
            .O(N__19445),
            .I(N__19437));
    LocalMux I__1884 (
            .O(N__19442),
            .I(N__19437));
    Span4Mux_v I__1883 (
            .O(N__19437),
            .I(N__19434));
    Odrv4 I__1882 (
            .O(N__19434),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    CascadeMux I__1881 (
            .O(N__19431),
            .I(N__19428));
    InMux I__1880 (
            .O(N__19428),
            .I(N__19425));
    LocalMux I__1879 (
            .O(N__19425),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__1878 (
            .O(N__19422),
            .I(N__19419));
    LocalMux I__1877 (
            .O(N__19419),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    CascadeMux I__1876 (
            .O(N__19416),
            .I(N__19413));
    InMux I__1875 (
            .O(N__19413),
            .I(N__19410));
    LocalMux I__1874 (
            .O(N__19410),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    CascadeMux I__1873 (
            .O(N__19407),
            .I(N__19404));
    InMux I__1872 (
            .O(N__19404),
            .I(N__19401));
    LocalMux I__1871 (
            .O(N__19401),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    CascadeMux I__1870 (
            .O(N__19398),
            .I(N__19395));
    InMux I__1869 (
            .O(N__19395),
            .I(N__19392));
    LocalMux I__1868 (
            .O(N__19392),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    CascadeMux I__1867 (
            .O(N__19389),
            .I(N__19386));
    InMux I__1866 (
            .O(N__19386),
            .I(N__19383));
    LocalMux I__1865 (
            .O(N__19383),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__1864 (
            .O(N__19380),
            .I(N__19377));
    InMux I__1863 (
            .O(N__19377),
            .I(N__19374));
    LocalMux I__1862 (
            .O(N__19374),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    CascadeMux I__1861 (
            .O(N__19371),
            .I(N__19367));
    CascadeMux I__1860 (
            .O(N__19370),
            .I(N__19364));
    InMux I__1859 (
            .O(N__19367),
            .I(N__19358));
    InMux I__1858 (
            .O(N__19364),
            .I(N__19358));
    CascadeMux I__1857 (
            .O(N__19363),
            .I(N__19355));
    LocalMux I__1856 (
            .O(N__19358),
            .I(N__19352));
    InMux I__1855 (
            .O(N__19355),
            .I(N__19349));
    Odrv4 I__1854 (
            .O(N__19352),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    LocalMux I__1853 (
            .O(N__19349),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1852 (
            .O(N__19344),
            .I(N__19340));
    InMux I__1851 (
            .O(N__19343),
            .I(N__19337));
    LocalMux I__1850 (
            .O(N__19340),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    LocalMux I__1849 (
            .O(N__19337),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    InMux I__1848 (
            .O(N__19332),
            .I(N__19320));
    InMux I__1847 (
            .O(N__19331),
            .I(N__19320));
    InMux I__1846 (
            .O(N__19330),
            .I(N__19320));
    InMux I__1845 (
            .O(N__19329),
            .I(N__19320));
    LocalMux I__1844 (
            .O(N__19320),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    CascadeMux I__1843 (
            .O(N__19317),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ));
    InMux I__1842 (
            .O(N__19314),
            .I(N__19311));
    LocalMux I__1841 (
            .O(N__19311),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    CascadeMux I__1840 (
            .O(N__19308),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ));
    InMux I__1839 (
            .O(N__19305),
            .I(N__19302));
    LocalMux I__1838 (
            .O(N__19302),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ));
    InMux I__1837 (
            .O(N__19299),
            .I(N__19296));
    LocalMux I__1836 (
            .O(N__19296),
            .I(N__19293));
    Odrv4 I__1835 (
            .O(N__19293),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ));
    CascadeMux I__1834 (
            .O(N__19290),
            .I(\current_shift_inst.PI_CTRL.N_98_cascade_ ));
    CascadeMux I__1833 (
            .O(N__19287),
            .I(\current_shift_inst.PI_CTRL.N_96_cascade_ ));
    InMux I__1832 (
            .O(N__19284),
            .I(N__19281));
    LocalMux I__1831 (
            .O(N__19281),
            .I(N__19278));
    Odrv12 I__1830 (
            .O(N__19278),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    CascadeMux I__1829 (
            .O(N__19275),
            .I(N__19272));
    InMux I__1828 (
            .O(N__19272),
            .I(N__19269));
    LocalMux I__1827 (
            .O(N__19269),
            .I(N__19266));
    Span4Mux_v I__1826 (
            .O(N__19266),
            .I(N__19263));
    Odrv4 I__1825 (
            .O(N__19263),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ));
    InMux I__1824 (
            .O(N__19260),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__1823 (
            .O(N__19257),
            .I(N__19254));
    LocalMux I__1822 (
            .O(N__19254),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__1821 (
            .O(N__19251),
            .I(N__19248));
    LocalMux I__1820 (
            .O(N__19248),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__1819 (
            .O(N__19245),
            .I(N__19242));
    InMux I__1818 (
            .O(N__19242),
            .I(N__19239));
    LocalMux I__1817 (
            .O(N__19239),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__1816 (
            .O(N__19236),
            .I(N__19233));
    LocalMux I__1815 (
            .O(N__19233),
            .I(N__19230));
    Odrv12 I__1814 (
            .O(N__19230),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    CascadeMux I__1813 (
            .O(N__19227),
            .I(N__19224));
    InMux I__1812 (
            .O(N__19224),
            .I(N__19221));
    LocalMux I__1811 (
            .O(N__19221),
            .I(N__19218));
    Odrv4 I__1810 (
            .O(N__19218),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    CascadeMux I__1809 (
            .O(N__19215),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ));
    InMux I__1808 (
            .O(N__19212),
            .I(N__19209));
    LocalMux I__1807 (
            .O(N__19209),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    CascadeMux I__1806 (
            .O(N__19206),
            .I(N__19203));
    InMux I__1805 (
            .O(N__19203),
            .I(N__19200));
    LocalMux I__1804 (
            .O(N__19200),
            .I(N__19197));
    Odrv12 I__1803 (
            .O(N__19197),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__1802 (
            .O(N__19194),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    InMux I__1801 (
            .O(N__19191),
            .I(N__19188));
    LocalMux I__1800 (
            .O(N__19188),
            .I(N__19185));
    Odrv12 I__1799 (
            .O(N__19185),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__1798 (
            .O(N__19182),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__1797 (
            .O(N__19179),
            .I(N__19176));
    InMux I__1796 (
            .O(N__19176),
            .I(N__19173));
    LocalMux I__1795 (
            .O(N__19173),
            .I(N__19170));
    Span4Mux_v I__1794 (
            .O(N__19170),
            .I(N__19167));
    Odrv4 I__1793 (
            .O(N__19167),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__1792 (
            .O(N__19164),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    CascadeMux I__1791 (
            .O(N__19161),
            .I(N__19158));
    InMux I__1790 (
            .O(N__19158),
            .I(N__19155));
    LocalMux I__1789 (
            .O(N__19155),
            .I(N__19152));
    Span4Mux_v I__1788 (
            .O(N__19152),
            .I(N__19149));
    Odrv4 I__1787 (
            .O(N__19149),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__1786 (
            .O(N__19146),
            .I(bfn_1_15_0_));
    CascadeMux I__1785 (
            .O(N__19143),
            .I(N__19140));
    InMux I__1784 (
            .O(N__19140),
            .I(N__19137));
    LocalMux I__1783 (
            .O(N__19137),
            .I(N__19134));
    Odrv12 I__1782 (
            .O(N__19134),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__1781 (
            .O(N__19131),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    CascadeMux I__1780 (
            .O(N__19128),
            .I(N__19125));
    InMux I__1779 (
            .O(N__19125),
            .I(N__19122));
    LocalMux I__1778 (
            .O(N__19122),
            .I(N__19119));
    Span4Mux_v I__1777 (
            .O(N__19119),
            .I(N__19116));
    Odrv4 I__1776 (
            .O(N__19116),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__1775 (
            .O(N__19113),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    CascadeMux I__1774 (
            .O(N__19110),
            .I(N__19107));
    InMux I__1773 (
            .O(N__19107),
            .I(N__19104));
    LocalMux I__1772 (
            .O(N__19104),
            .I(N__19101));
    Odrv12 I__1771 (
            .O(N__19101),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__1770 (
            .O(N__19098),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    InMux I__1769 (
            .O(N__19095),
            .I(N__19092));
    LocalMux I__1768 (
            .O(N__19092),
            .I(N__19089));
    Odrv12 I__1767 (
            .O(N__19089),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__1766 (
            .O(N__19086),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__1765 (
            .O(N__19083),
            .I(N__19080));
    InMux I__1764 (
            .O(N__19080),
            .I(N__19077));
    LocalMux I__1763 (
            .O(N__19077),
            .I(N__19074));
    Span4Mux_v I__1762 (
            .O(N__19074),
            .I(N__19071));
    Odrv4 I__1761 (
            .O(N__19071),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__1760 (
            .O(N__19068),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    CascadeMux I__1759 (
            .O(N__19065),
            .I(N__19062));
    InMux I__1758 (
            .O(N__19062),
            .I(N__19059));
    LocalMux I__1757 (
            .O(N__19059),
            .I(N__19056));
    Odrv4 I__1756 (
            .O(N__19056),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__1755 (
            .O(N__19053),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__1754 (
            .O(N__19050),
            .I(N__19047));
    InMux I__1753 (
            .O(N__19047),
            .I(N__19044));
    LocalMux I__1752 (
            .O(N__19044),
            .I(N__19041));
    Odrv4 I__1751 (
            .O(N__19041),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__1750 (
            .O(N__19038),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__1749 (
            .O(N__19035),
            .I(N__19032));
    InMux I__1748 (
            .O(N__19032),
            .I(N__19029));
    LocalMux I__1747 (
            .O(N__19029),
            .I(N__19026));
    Span4Mux_v I__1746 (
            .O(N__19026),
            .I(N__19023));
    Odrv4 I__1745 (
            .O(N__19023),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__1744 (
            .O(N__19020),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    CascadeMux I__1743 (
            .O(N__19017),
            .I(N__19014));
    InMux I__1742 (
            .O(N__19014),
            .I(N__19011));
    LocalMux I__1741 (
            .O(N__19011),
            .I(N__19008));
    Span4Mux_v I__1740 (
            .O(N__19008),
            .I(N__19005));
    Odrv4 I__1739 (
            .O(N__19005),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__1738 (
            .O(N__19002),
            .I(bfn_1_14_0_));
    InMux I__1737 (
            .O(N__18999),
            .I(N__18996));
    LocalMux I__1736 (
            .O(N__18996),
            .I(N__18993));
    Odrv12 I__1735 (
            .O(N__18993),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__1734 (
            .O(N__18990),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__1733 (
            .O(N__18987),
            .I(N__18984));
    InMux I__1732 (
            .O(N__18984),
            .I(N__18981));
    LocalMux I__1731 (
            .O(N__18981),
            .I(N__18978));
    Odrv12 I__1730 (
            .O(N__18978),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__1729 (
            .O(N__18975),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    CascadeMux I__1728 (
            .O(N__18972),
            .I(N__18969));
    InMux I__1727 (
            .O(N__18969),
            .I(N__18966));
    LocalMux I__1726 (
            .O(N__18966),
            .I(N__18963));
    Odrv12 I__1725 (
            .O(N__18963),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__1724 (
            .O(N__18960),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__1723 (
            .O(N__18957),
            .I(N__18954));
    InMux I__1722 (
            .O(N__18954),
            .I(N__18951));
    LocalMux I__1721 (
            .O(N__18951),
            .I(N__18948));
    Odrv12 I__1720 (
            .O(N__18948),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__1719 (
            .O(N__18945),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    InMux I__1718 (
            .O(N__18942),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__1717 (
            .O(N__18939),
            .I(N__18936));
    InMux I__1716 (
            .O(N__18936),
            .I(N__18933));
    LocalMux I__1715 (
            .O(N__18933),
            .I(N__18930));
    Odrv4 I__1714 (
            .O(N__18930),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__1713 (
            .O(N__18927),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__1712 (
            .O(N__18924),
            .I(N__18921));
    InMux I__1711 (
            .O(N__18921),
            .I(N__18918));
    LocalMux I__1710 (
            .O(N__18918),
            .I(N__18915));
    Span4Mux_h I__1709 (
            .O(N__18915),
            .I(N__18912));
    Odrv4 I__1708 (
            .O(N__18912),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__1707 (
            .O(N__18909),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__1706 (
            .O(N__18906),
            .I(N__18903));
    InMux I__1705 (
            .O(N__18903),
            .I(N__18900));
    LocalMux I__1704 (
            .O(N__18900),
            .I(N__18897));
    Span4Mux_v I__1703 (
            .O(N__18897),
            .I(N__18894));
    Odrv4 I__1702 (
            .O(N__18894),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__1701 (
            .O(N__18891),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    InMux I__1700 (
            .O(N__18888),
            .I(N__18885));
    LocalMux I__1699 (
            .O(N__18885),
            .I(N__18882));
    Span4Mux_h I__1698 (
            .O(N__18882),
            .I(N__18879));
    Odrv4 I__1697 (
            .O(N__18879),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    InMux I__1696 (
            .O(N__18876),
            .I(bfn_1_13_0_));
    CascadeMux I__1695 (
            .O(N__18873),
            .I(N__18870));
    InMux I__1694 (
            .O(N__18870),
            .I(N__18867));
    LocalMux I__1693 (
            .O(N__18867),
            .I(N__18864));
    Span4Mux_h I__1692 (
            .O(N__18864),
            .I(N__18861));
    Odrv4 I__1691 (
            .O(N__18861),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__1690 (
            .O(N__18858),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__1689 (
            .O(N__18855),
            .I(N__18852));
    InMux I__1688 (
            .O(N__18852),
            .I(N__18849));
    LocalMux I__1687 (
            .O(N__18849),
            .I(N__18846));
    Span4Mux_v I__1686 (
            .O(N__18846),
            .I(N__18843));
    Span4Mux_s1_h I__1685 (
            .O(N__18843),
            .I(N__18840));
    Odrv4 I__1684 (
            .O(N__18840),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__1683 (
            .O(N__18837),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    CascadeMux I__1682 (
            .O(N__18834),
            .I(N__18831));
    InMux I__1681 (
            .O(N__18831),
            .I(N__18828));
    LocalMux I__1680 (
            .O(N__18828),
            .I(N__18825));
    Span4Mux_v I__1679 (
            .O(N__18825),
            .I(N__18822));
    Odrv4 I__1678 (
            .O(N__18822),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__1677 (
            .O(N__18819),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__1676 (
            .O(N__18816),
            .I(N__18813));
    InMux I__1675 (
            .O(N__18813),
            .I(N__18810));
    LocalMux I__1674 (
            .O(N__18810),
            .I(N__18807));
    Odrv4 I__1673 (
            .O(N__18807),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__1672 (
            .O(N__18804),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    InMux I__1671 (
            .O(N__18801),
            .I(N__18798));
    LocalMux I__1670 (
            .O(N__18798),
            .I(N__18795));
    Span4Mux_v I__1669 (
            .O(N__18795),
            .I(N__18792));
    Odrv4 I__1668 (
            .O(N__18792),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    InMux I__1667 (
            .O(N__18789),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__1666 (
            .O(N__18786),
            .I(N__18783));
    LocalMux I__1665 (
            .O(N__18783),
            .I(N__18780));
    Span4Mux_v I__1664 (
            .O(N__18780),
            .I(N__18777));
    Odrv4 I__1663 (
            .O(N__18777),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    InMux I__1662 (
            .O(N__18774),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    InMux I__1661 (
            .O(N__18771),
            .I(N__18768));
    LocalMux I__1660 (
            .O(N__18768),
            .I(N__18765));
    Span4Mux_v I__1659 (
            .O(N__18765),
            .I(N__18762));
    Odrv4 I__1658 (
            .O(N__18762),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    CascadeMux I__1657 (
            .O(N__18759),
            .I(N__18754));
    CascadeMux I__1656 (
            .O(N__18758),
            .I(N__18750));
    InMux I__1655 (
            .O(N__18757),
            .I(N__18741));
    InMux I__1654 (
            .O(N__18754),
            .I(N__18741));
    InMux I__1653 (
            .O(N__18753),
            .I(N__18741));
    InMux I__1652 (
            .O(N__18750),
            .I(N__18741));
    LocalMux I__1651 (
            .O(N__18741),
            .I(N__18730));
    CascadeMux I__1650 (
            .O(N__18740),
            .I(N__18727));
    CascadeMux I__1649 (
            .O(N__18739),
            .I(N__18724));
    CascadeMux I__1648 (
            .O(N__18738),
            .I(N__18721));
    CascadeMux I__1647 (
            .O(N__18737),
            .I(N__18718));
    CascadeMux I__1646 (
            .O(N__18736),
            .I(N__18715));
    CascadeMux I__1645 (
            .O(N__18735),
            .I(N__18712));
    CascadeMux I__1644 (
            .O(N__18734),
            .I(N__18709));
    InMux I__1643 (
            .O(N__18733),
            .I(N__18706));
    Span4Mux_v I__1642 (
            .O(N__18730),
            .I(N__18703));
    InMux I__1641 (
            .O(N__18727),
            .I(N__18696));
    InMux I__1640 (
            .O(N__18724),
            .I(N__18696));
    InMux I__1639 (
            .O(N__18721),
            .I(N__18696));
    InMux I__1638 (
            .O(N__18718),
            .I(N__18687));
    InMux I__1637 (
            .O(N__18715),
            .I(N__18687));
    InMux I__1636 (
            .O(N__18712),
            .I(N__18687));
    InMux I__1635 (
            .O(N__18709),
            .I(N__18687));
    LocalMux I__1634 (
            .O(N__18706),
            .I(N__18682));
    Span4Mux_s1_h I__1633 (
            .O(N__18703),
            .I(N__18682));
    LocalMux I__1632 (
            .O(N__18696),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1631 (
            .O(N__18687),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    Odrv4 I__1630 (
            .O(N__18682),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    InMux I__1629 (
            .O(N__18675),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__1628 (
            .O(N__18672),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    CascadeMux I__1627 (
            .O(N__18669),
            .I(N__18666));
    InMux I__1626 (
            .O(N__18666),
            .I(N__18663));
    LocalMux I__1625 (
            .O(N__18663),
            .I(N__18660));
    Span4Mux_v I__1624 (
            .O(N__18660),
            .I(N__18657));
    Odrv4 I__1623 (
            .O(N__18657),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__1622 (
            .O(N__18654),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    InMux I__1621 (
            .O(N__18651),
            .I(N__18648));
    LocalMux I__1620 (
            .O(N__18648),
            .I(N__18645));
    Odrv4 I__1619 (
            .O(N__18645),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__1618 (
            .O(N__18642),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__1617 (
            .O(N__18639),
            .I(N__18636));
    InMux I__1616 (
            .O(N__18636),
            .I(N__18633));
    LocalMux I__1615 (
            .O(N__18633),
            .I(N__18630));
    Odrv4 I__1614 (
            .O(N__18630),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    InMux I__1613 (
            .O(N__18627),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    CascadeMux I__1612 (
            .O(N__18624),
            .I(N__18621));
    InMux I__1611 (
            .O(N__18621),
            .I(N__18618));
    LocalMux I__1610 (
            .O(N__18618),
            .I(N__18615));
    Span4Mux_h I__1609 (
            .O(N__18615),
            .I(N__18612));
    Odrv4 I__1608 (
            .O(N__18612),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__1607 (
            .O(N__18609),
            .I(N__18606));
    LocalMux I__1606 (
            .O(N__18606),
            .I(N__18603));
    Span4Mux_v I__1605 (
            .O(N__18603),
            .I(N__18600));
    Odrv4 I__1604 (
            .O(N__18600),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    InMux I__1603 (
            .O(N__18597),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    CascadeMux I__1602 (
            .O(N__18594),
            .I(N__18591));
    InMux I__1601 (
            .O(N__18591),
            .I(N__18588));
    LocalMux I__1600 (
            .O(N__18588),
            .I(N__18585));
    Span4Mux_v I__1599 (
            .O(N__18585),
            .I(N__18582));
    Odrv4 I__1598 (
            .O(N__18582),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    InMux I__1597 (
            .O(N__18579),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__1596 (
            .O(N__18576),
            .I(N__18573));
    LocalMux I__1595 (
            .O(N__18573),
            .I(N__18570));
    Span4Mux_v I__1594 (
            .O(N__18570),
            .I(N__18567));
    Odrv4 I__1593 (
            .O(N__18567),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    InMux I__1592 (
            .O(N__18564),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    CascadeMux I__1591 (
            .O(N__18561),
            .I(N__18558));
    InMux I__1590 (
            .O(N__18558),
            .I(N__18555));
    LocalMux I__1589 (
            .O(N__18555),
            .I(N__18552));
    Span4Mux_v I__1588 (
            .O(N__18552),
            .I(N__18549));
    Odrv4 I__1587 (
            .O(N__18549),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__1586 (
            .O(N__18546),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    InMux I__1585 (
            .O(N__18543),
            .I(N__18540));
    LocalMux I__1584 (
            .O(N__18540),
            .I(N__18537));
    Span4Mux_v I__1583 (
            .O(N__18537),
            .I(N__18534));
    Odrv4 I__1582 (
            .O(N__18534),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    InMux I__1581 (
            .O(N__18531),
            .I(bfn_1_11_0_));
    InMux I__1580 (
            .O(N__18528),
            .I(N__18525));
    LocalMux I__1579 (
            .O(N__18525),
            .I(N__18522));
    Span4Mux_v I__1578 (
            .O(N__18522),
            .I(N__18519));
    Odrv4 I__1577 (
            .O(N__18519),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    InMux I__1576 (
            .O(N__18516),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    InMux I__1575 (
            .O(N__18513),
            .I(N__18510));
    LocalMux I__1574 (
            .O(N__18510),
            .I(N__18507));
    Span4Mux_v I__1573 (
            .O(N__18507),
            .I(N__18504));
    Span4Mux_s1_h I__1572 (
            .O(N__18504),
            .I(N__18501));
    Odrv4 I__1571 (
            .O(N__18501),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__1570 (
            .O(N__18498),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__1569 (
            .O(N__18495),
            .I(N__18492));
    LocalMux I__1568 (
            .O(N__18492),
            .I(N__18489));
    Span4Mux_v I__1567 (
            .O(N__18489),
            .I(N__18486));
    Odrv4 I__1566 (
            .O(N__18486),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__1565 (
            .O(N__18483),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__1564 (
            .O(N__18480),
            .I(N__18477));
    LocalMux I__1563 (
            .O(N__18477),
            .I(N__18474));
    Odrv4 I__1562 (
            .O(N__18474),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    InMux I__1561 (
            .O(N__18471),
            .I(N__18468));
    LocalMux I__1560 (
            .O(N__18468),
            .I(N__18465));
    Span4Mux_v I__1559 (
            .O(N__18465),
            .I(N__18462));
    Odrv4 I__1558 (
            .O(N__18462),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__1557 (
            .O(N__18459),
            .I(N__18456));
    InMux I__1556 (
            .O(N__18456),
            .I(N__18453));
    LocalMux I__1555 (
            .O(N__18453),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    InMux I__1554 (
            .O(N__18450),
            .I(N__18447));
    LocalMux I__1553 (
            .O(N__18447),
            .I(N__18444));
    Span4Mux_v I__1552 (
            .O(N__18444),
            .I(N__18441));
    Odrv4 I__1551 (
            .O(N__18441),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__1550 (
            .O(N__18438),
            .I(N__18435));
    InMux I__1549 (
            .O(N__18435),
            .I(N__18432));
    LocalMux I__1548 (
            .O(N__18432),
            .I(N__18429));
    Odrv4 I__1547 (
            .O(N__18429),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    InMux I__1546 (
            .O(N__18426),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__1545 (
            .O(N__18423),
            .I(N__18420));
    LocalMux I__1544 (
            .O(N__18420),
            .I(N__18417));
    Span4Mux_v I__1543 (
            .O(N__18417),
            .I(N__18414));
    Odrv4 I__1542 (
            .O(N__18414),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__1541 (
            .O(N__18411),
            .I(N__18408));
    InMux I__1540 (
            .O(N__18408),
            .I(N__18405));
    LocalMux I__1539 (
            .O(N__18405),
            .I(N__18402));
    Odrv4 I__1538 (
            .O(N__18402),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    InMux I__1537 (
            .O(N__18399),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    InMux I__1536 (
            .O(N__18396),
            .I(N__18393));
    LocalMux I__1535 (
            .O(N__18393),
            .I(N__18390));
    Span4Mux_v I__1534 (
            .O(N__18390),
            .I(N__18387));
    Odrv4 I__1533 (
            .O(N__18387),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__1532 (
            .O(N__18384),
            .I(N__18381));
    InMux I__1531 (
            .O(N__18381),
            .I(N__18378));
    LocalMux I__1530 (
            .O(N__18378),
            .I(N__18375));
    Odrv4 I__1529 (
            .O(N__18375),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__1528 (
            .O(N__18372),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    IoInMux I__1527 (
            .O(N__18369),
            .I(N__18366));
    LocalMux I__1526 (
            .O(N__18366),
            .I(N__18363));
    Span4Mux_s3_v I__1525 (
            .O(N__18363),
            .I(N__18360));
    Span4Mux_h I__1524 (
            .O(N__18360),
            .I(N__18357));
    Sp12to4 I__1523 (
            .O(N__18357),
            .I(N__18354));
    Span12Mux_s9_v I__1522 (
            .O(N__18354),
            .I(N__18351));
    Span12Mux_v I__1521 (
            .O(N__18351),
            .I(N__18348));
    Odrv12 I__1520 (
            .O(N__18348),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1519 (
            .O(N__18345),
            .I(N__18342));
    LocalMux I__1518 (
            .O(N__18342),
            .I(N__18339));
    IoSpan4Mux I__1517 (
            .O(N__18339),
            .I(N__18336));
    IoSpan4Mux I__1516 (
            .O(N__18336),
            .I(N__18333));
    Odrv4 I__1515 (
            .O(N__18333),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_9_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_26_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_10_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_26_0_));
    defparam IN_MUX_bfv_10_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_27_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_10_27_0_));
    defparam IN_MUX_bfv_10_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_28_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_10_28_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_11_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_25_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_11_25_0_));
    defparam IN_MUX_bfv_7_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_26_0_));
    defparam IN_MUX_bfv_7_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_27_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_7_27_0_));
    defparam IN_MUX_bfv_7_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_28_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_7_28_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_17_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_17_22_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_5_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_5_16_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18369),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18345),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__33000),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_162_i_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__42123),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un1_start_g ));
    ICE_GB \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0  (
            .USERSIGNALTOGLOBALBUFFER(N__32487),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_hc.un1_start_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__35640),
            .CLKHFEN(N__35642),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__35641),
            .RGB2PWM(N__19461),
            .RGB1(rgb_g),
            .CURREN(N__35675),
            .RGB2(rgb_b),
            .RGB1PWM(N__20028),
            .RGB0PWM(N__47124),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(N__18480),
            .in2(_gnd_net_),
            .in3(N__18733),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__18471),
            .in2(N__18459),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__18450),
            .in2(N__18438),
            .in3(N__18426),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__18423),
            .in2(N__18411),
            .in3(N__18399),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__18396),
            .in2(N__18384),
            .in3(N__18372),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__18609),
            .in2(N__18758),
            .in3(N__18597),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__18753),
            .in2(N__18594),
            .in3(N__18579),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__18576),
            .in2(N__18759),
            .in3(N__18564),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__18757),
            .in2(N__18561),
            .in3(N__18546),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__18543),
            .in2(N__18734),
            .in3(N__18531),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__18528),
            .in2(N__18738),
            .in3(N__18516),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__18513),
            .in2(N__18735),
            .in3(N__18498),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__18495),
            .in2(N__18739),
            .in3(N__18483),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__18801),
            .in2(N__18736),
            .in3(N__18789),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__18786),
            .in2(N__18740),
            .in3(N__18774),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__18771),
            .in2(N__18737),
            .in3(N__18675),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18672),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__20187),
            .in2(N__19454),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__20155),
            .in2(N__18669),
            .in3(N__18654),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__18651),
            .in2(N__21094),
            .in3(N__18642),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__21022),
            .in2(N__18639),
            .in3(N__18627),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__20942),
            .in2(N__18624),
            .in3(N__18942),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__20862),
            .in2(N__18939),
            .in3(N__18927),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__20795),
            .in2(N__18924),
            .in3(N__18909),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(N__20727),
            .in2(N__18906),
            .in3(N__18891),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__18888),
            .in2(N__20654),
            .in3(N__18876),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__21529),
            .in2(N__18873),
            .in3(N__18858),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__21477),
            .in2(N__18855),
            .in3(N__18837),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__21436),
            .in2(N__18834),
            .in3(N__18819),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__21370),
            .in2(N__18816),
            .in3(N__18804),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__21308),
            .in2(N__19065),
            .in3(N__19053),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__21247),
            .in2(N__19050),
            .in3(N__19038),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__21195),
            .in2(N__19035),
            .in3(N__19020),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__21141),
            .in2(N__19017),
            .in3(N__19002),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__18999),
            .in2(N__21860),
            .in3(N__18990),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__21804),
            .in2(N__18987),
            .in3(N__18975),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__22773),
            .in2(N__18972),
            .in3(N__18960),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__22744),
            .in2(N__18957),
            .in3(N__18945),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__21768),
            .in2(N__19206),
            .in3(N__19194),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__19191),
            .in2(N__21720),
            .in3(N__19182),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__22815),
            .in2(N__19179),
            .in3(N__19164),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__21639),
            .in2(N__19161),
            .in3(N__19146),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__21591),
            .in2(N__19143),
            .in3(N__19131),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__22110),
            .in2(N__19128),
            .in3(N__19113),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__22071),
            .in2(N__19110),
            .in3(N__19098),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__19095),
            .in2(N__22030),
            .in3(N__19086),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__21982),
            .in2(N__19083),
            .in3(N__19068),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6  (
            .in0(N__19284),
            .in1(N__22620),
            .in2(N__19275),
            .in3(N__19260),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_0 .LUT_INIT=16'b1101110111001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_0  (
            .in0(N__20551),
            .in1(N__19257),
            .in2(N__20368),
            .in3(N__22652),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47516),
            .ce(),
            .sr(N__47089));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_2 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_2  (
            .in0(N__20552),
            .in1(N__22650),
            .in2(N__20369),
            .in3(N__19251),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47516),
            .ce(),
            .sr(N__47089));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5  (
            .in0(N__22649),
            .in1(N__20555),
            .in2(N__19245),
            .in3(N__20315),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47516),
            .ce(),
            .sr(N__47089));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_1_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_1_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_1_16_6 .LUT_INIT=16'b1011101100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_1_16_6  (
            .in0(N__20553),
            .in1(N__22651),
            .in2(N__20370),
            .in3(N__19236),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47516),
            .ce(),
            .sr(N__47089));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_1_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_1_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_1_16_7 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_1_16_7  (
            .in0(N__22648),
            .in1(N__20554),
            .in2(N__19227),
            .in3(N__20314),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47516),
            .ce(),
            .sr(N__47089));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_1_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_1_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_1_17_0  (
            .in0(N__21251),
            .in1(N__21371),
            .in2(N__21551),
            .in3(N__22034),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_1_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_1_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_1_17_1  (
            .in0(N__19212),
            .in1(N__19551),
            .in2(N__19215),
            .in3(N__19314),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_1_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_1_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_1_17_2  (
            .in0(N__21209),
            .in1(N__21309),
            .in2(N__21441),
            .in3(N__21494),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_1_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_1_18_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_1_18_2  (
            .in0(N__21858),
            .in1(N__21817),
            .in2(N__21161),
            .in3(N__21773),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_1_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_1_18_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_1_18_3  (
            .in0(N__22664),
            .in1(N__21724),
            .in2(N__19317),
            .in3(N__19299),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_1_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_1_19_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__21592),
            .in2(_gnd_net_),
            .in3(N__22737),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_1_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_1_19_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_1_19_2  (
            .in0(N__22076),
            .in1(N__22121),
            .in2(N__21651),
            .in3(N__21986),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_1_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_1_19_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_1_19_3  (
            .in0(N__22831),
            .in1(N__22786),
            .in2(N__19308),
            .in3(N__19305),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_1_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_1_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_1_21_1 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_1_21_1  (
            .in0(N__26902),
            .in1(N__20995),
            .in2(_gnd_net_),
            .in3(N__19907),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_5  (
            .in0(_gnd_net_),
            .in1(N__20994),
            .in2(_gnd_net_),
            .in3(N__21064),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_6 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_6  (
            .in0(N__19886),
            .in1(N__26903),
            .in2(N__19290),
            .in3(N__19677),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(\current_shift_inst.PI_CTRL.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_21_7 .LUT_INIT=16'b0000000011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_21_7  (
            .in0(N__19343),
            .in1(N__19946),
            .in2(N__19287),
            .in3(N__21065),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_0 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_0  (
            .in0(N__19639),
            .in1(N__21951),
            .in2(N__19370),
            .in3(N__19330),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__47098));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_1 .LUT_INIT=16'b1111010101000100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_1  (
            .in0(N__26908),
            .in1(N__19960),
            .in2(N__19701),
            .in3(N__20931),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__47098));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_2 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_2  (
            .in0(N__19640),
            .in1(N__20583),
            .in2(N__19371),
            .in3(N__19331),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__47098));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3  (
            .in0(N__19329),
            .in1(N__20130),
            .in2(N__19363),
            .in3(N__19641),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__47098));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4 .LUT_INIT=16'b1010101011111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4  (
            .in0(N__21069),
            .in1(N__19344),
            .in2(N__19965),
            .in3(N__19332),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__47098));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6  (
            .in0(N__21003),
            .in1(N__19896),
            .in2(N__19702),
            .in3(N__19887),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__47098));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_0 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_0  (
            .in0(N__26909),
            .in1(N__20844),
            .in2(N__19703),
            .in3(N__19963),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47442),
            .ce(),
            .sr(N__47099));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_1 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_1  (
            .in0(N__19961),
            .in1(N__26910),
            .in2(N__20769),
            .in3(N__19699),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47442),
            .ce(),
            .sr(N__47099));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_2 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_2  (
            .in0(N__26911),
            .in1(N__20691),
            .in2(N__19704),
            .in3(N__19964),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47442),
            .ce(),
            .sr(N__47099));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_7 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_7  (
            .in0(N__19962),
            .in1(N__26912),
            .in2(N__20622),
            .in3(N__19700),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47442),
            .ce(),
            .sr(N__47099));
    defparam rgb_drv_RNO_0_LC_1_30_6.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_1_30_6.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_1_30_6.LUT_INIT=16'b1010101001010101;
    LogicCell40 rgb_drv_RNO_0_LC_1_30_6 (
            .in0(N__47123),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32673),
            .lcout(N_38_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_6 .LUT_INIT=16'b0101101001001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_6  (
            .in0(N__20194),
            .in1(N__20523),
            .in2(N__19455),
            .in3(N__20378),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47547),
            .ce(),
            .sr(N__47071));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_0 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_0  (
            .in0(N__22691),
            .in1(N__20520),
            .in2(N__19431),
            .in3(N__20375),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47538),
            .ce(),
            .sr(N__47074));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_1  (
            .in0(N__20518),
            .in1(N__20371),
            .in2(_gnd_net_),
            .in3(N__19422),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47538),
            .ce(),
            .sr(N__47074));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_2_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_2_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_2_13_3 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_2_13_3  (
            .in0(N__20516),
            .in1(N__22694),
            .in2(N__19416),
            .in3(N__20372),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47538),
            .ce(),
            .sr(N__47074));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_2_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_2_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_2_13_4 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_2_13_4  (
            .in0(N__22692),
            .in1(N__20521),
            .in2(N__19407),
            .in3(N__20376),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47538),
            .ce(),
            .sr(N__47074));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_5 .LUT_INIT=16'b1011000010110001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_5  (
            .in0(N__20519),
            .in1(N__22696),
            .in2(N__19398),
            .in3(N__20374),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47538),
            .ce(),
            .sr(N__47074));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_2_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_2_13_6 .LUT_INIT=16'b1101000011010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_2_13_6  (
            .in0(N__22693),
            .in1(N__20522),
            .in2(N__19389),
            .in3(N__20377),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47538),
            .ce(),
            .sr(N__47074));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_7 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_7  (
            .in0(N__20517),
            .in1(N__22695),
            .in2(N__19380),
            .in3(N__20373),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47538),
            .ce(),
            .sr(N__47074));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_0 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_0  (
            .in0(N__22699),
            .in1(N__20514),
            .in2(N__20399),
            .in3(N__19539),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47529),
            .ce(),
            .sr(N__47079));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1  (
            .in0(N__20512),
            .in1(N__22702),
            .in2(N__19533),
            .in3(N__20395),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47529),
            .ce(),
            .sr(N__47079));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_2 .LUT_INIT=16'b1100110011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_2  (
            .in0(N__22700),
            .in1(N__19524),
            .in2(N__20400),
            .in3(N__20515),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47529),
            .ce(),
            .sr(N__47079));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_5 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_5  (
            .in0(N__20511),
            .in1(N__22701),
            .in2(N__19515),
            .in3(N__20394),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47529),
            .ce(),
            .sr(N__47079));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_7 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_7  (
            .in0(N__20513),
            .in1(N__22703),
            .in2(N__19506),
            .in3(N__20396),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47529),
            .ce(),
            .sr(N__47079));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_0 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_0  (
            .in0(N__22655),
            .in1(N__20525),
            .in2(N__19494),
            .in3(N__20355),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47517),
            .ce(),
            .sr(N__47083));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_2_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_2_15_1 .LUT_INIT=16'b1111001111100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_2_15_1  (
            .in0(N__20350),
            .in1(N__20557),
            .in2(N__19485),
            .in3(N__22660),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47517),
            .ce(),
            .sr(N__47083));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_2_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_2_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_2_15_2 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_2_15_2  (
            .in0(N__22656),
            .in1(N__20526),
            .in2(N__19476),
            .in3(N__20356),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47517),
            .ce(),
            .sr(N__47083));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_3 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_3  (
            .in0(N__20351),
            .in1(N__22657),
            .in2(N__20558),
            .in3(N__19467),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47517),
            .ce(),
            .sr(N__47083));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_5 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_5  (
            .in0(N__20352),
            .in1(N__22658),
            .in2(N__20559),
            .in3(N__19593),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47517),
            .ce(),
            .sr(N__47083));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_6 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_6  (
            .in0(N__22654),
            .in1(N__20524),
            .in2(N__19587),
            .in3(N__20354),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47517),
            .ce(),
            .sr(N__47083));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_7 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_7  (
            .in0(N__20353),
            .in1(N__22659),
            .in2(N__20560),
            .in3(N__19578),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47517),
            .ce(),
            .sr(N__47083));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_2_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_2_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_2_16_2 .LUT_INIT=16'b1101000011010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_2_16_2  (
            .in0(N__22653),
            .in1(N__20556),
            .in2(N__19572),
            .in3(N__20316),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47504),
            .ce(),
            .sr(N__47087));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__21300),
            .in2(_gnd_net_),
            .in3(N__21487),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_2_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_2_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_2_17_1  (
            .in0(N__21437),
            .in1(N__19608),
            .in2(N__19557),
            .in3(N__21981),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_17_3 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_17_3  (
            .in0(N__21106),
            .in1(N__20165),
            .in2(N__20209),
            .in3(N__21034),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_4 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_4  (
            .in0(N__19545),
            .in1(N__20647),
            .in2(N__19554),
            .in3(N__20878),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5  (
            .in0(N__20790),
            .in1(N__20956),
            .in2(_gnd_net_),
            .in3(N__20728),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_2_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_2_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_2_17_6  (
            .in0(N__20729),
            .in1(N__20791),
            .in2(N__20882),
            .in3(N__20646),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_17_7 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_17_7  (
            .in0(N__21107),
            .in1(N__21035),
            .in2(N__19629),
            .in3(N__20957),
            .lcout(\current_shift_inst.PI_CTRL.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_18_3  (
            .in0(N__21769),
            .in1(N__21859),
            .in2(N__21824),
            .in3(N__21160),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_18_4  (
            .in0(N__22026),
            .in1(N__21731),
            .in2(N__19626),
            .in3(N__19623),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_2_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_2_18_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_2_18_5  (
            .in0(N__19617),
            .in1(N__22554),
            .in2(N__19611),
            .in3(N__19602),
            .lcout(\current_shift_inst.PI_CTRL.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_2_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_2_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_2_18_6  (
            .in0(N__21243),
            .in1(N__21360),
            .in2(N__21210),
            .in3(N__21535),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_2_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_2_18_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_2_18_7  (
            .in0(N__22117),
            .in1(N__21643),
            .in2(N__21608),
            .in3(N__22072),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_3  (
            .in0(N__21326),
            .in1(N__21668),
            .in2(N__21687),
            .in3(N__21272),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_20_0 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_20_0  (
            .in0(N__20608),
            .in1(_gnd_net_),
            .in2(N__20926),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_1  (
            .in0(N__20683),
            .in1(N__20764),
            .in2(N__19596),
            .in3(N__20833),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_20_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(N__21398),
            .in2(_gnd_net_),
            .in3(N__21887),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_20_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_20_4  (
            .in0(N__21458),
            .in1(N__22326),
            .in2(N__19728),
            .in3(N__19725),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_20_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_20_5  (
            .in0(N__21273),
            .in1(N__21935),
            .in2(N__21330),
            .in3(N__21920),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_20_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_20_6  (
            .in0(N__21669),
            .in1(N__21683),
            .in2(N__22343),
            .in3(N__21902),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_0  (
            .in0(N__22242),
            .in1(N__19719),
            .in2(N__19713),
            .in3(N__22371),
            .lcout(\current_shift_inst.PI_CTRL.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_21_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_21_5  (
            .in0(_gnd_net_),
            .in1(N__22404),
            .in2(_gnd_net_),
            .in3(N__22389),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_21_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_21_6  (
            .in0(N__21459),
            .in1(N__21402),
            .in2(N__19656),
            .in3(N__21870),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_21_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_21_7  (
            .in0(N__21909),
            .in1(N__19653),
            .in2(N__19644),
            .in3(N__22308),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_3 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_3  (
            .in0(_gnd_net_),
            .in1(N__19913),
            .in2(N__26904),
            .in3(N__19945),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_22_4 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_22_4  (
            .in0(N__21002),
            .in1(N__19947),
            .in2(N__19917),
            .in3(N__26886),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_22_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_22_5  (
            .in0(_gnd_net_),
            .in1(N__20687),
            .in2(_gnd_net_),
            .in3(N__20927),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_22_6  (
            .in0(N__20765),
            .in1(N__20840),
            .in2(N__19890),
            .in3(N__20615),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_0  (
            .in0(N__19871),
            .in1(N__19856),
            .in2(_gnd_net_),
            .in3(N__19838),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3  (
            .in0(N__19753),
            .in1(N__19823),
            .in2(N__19784),
            .in3(N__19801),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_5  (
            .in0(_gnd_net_),
            .in1(N__19822),
            .in2(_gnd_net_),
            .in3(N__20047),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_6  (
            .in0(N__19802),
            .in1(N__19780),
            .in2(N__19761),
            .in3(N__19754),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_7 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_7  (
            .in0(N__19737),
            .in1(N__20074),
            .in2(N__19731),
            .in3(N__20101),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_24_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_24_5 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_24_5  (
            .in0(N__20112),
            .in1(N__20106),
            .in2(N__20082),
            .in3(N__20054),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_LC_2_30_2.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_2_30_2.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_2_30_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_drv_RNO_LC_2_30_2 (
            .in0(N__47122),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32672),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_4  (
            .in0(N__20019),
            .in1(N__20568),
            .in2(_gnd_net_),
            .in3(N__20397),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47539),
            .ce(),
            .sr(N__47067));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_13_7 .LUT_INIT=16'b1101000011010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_3_13_7  (
            .in0(N__22704),
            .in1(N__20561),
            .in2(N__20010),
            .in3(N__20398),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47530),
            .ce(),
            .sr(N__47072));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_3_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_3_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_3_14_2 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_3_14_2  (
            .in0(N__20386),
            .in1(N__22705),
            .in2(N__19995),
            .in3(N__20565),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47518),
            .ce(),
            .sr(N__47075));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_3_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_3_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_3_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22538),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47505),
            .ce(),
            .sr(N__47080));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23027),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47505),
            .ce(),
            .sr(N__47080));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_15_5 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_3_15_5  (
            .in0(N__22698),
            .in1(N__20567),
            .in2(N__19980),
            .in3(N__20385),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47505),
            .ce(),
            .sr(N__47080));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22490),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47505),
            .ce(),
            .sr(N__47080));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_3_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_3_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_3_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22433),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47492),
            .ce(),
            .sr(N__47084));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22949),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47492),
            .ce(),
            .sr(N__47084));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_3_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_3_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_3_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22922),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47492),
            .ce(),
            .sr(N__47084));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_3_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_3_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_3_16_3 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_3_16_3  (
            .in0(N__20228),
            .in1(N__20213),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47492),
            .ce(),
            .sr(N__47084));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_3_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_3_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_3_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_3_16_4  (
            .in0(N__22467),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47492),
            .ce(),
            .sr(N__47084));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_3_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_3_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_3_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22871),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47492),
            .ce(),
            .sr(N__47084));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_3_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_3_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_3_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23003),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47492),
            .ce(),
            .sr(N__47084));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_16_7 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_3_16_7  (
            .in0(N__22706),
            .in1(N__20566),
            .in2(N__20415),
            .in3(N__20387),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47492),
            .ce(),
            .sr(N__47084));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__20229),
            .in2(N__20214),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__22236),
            .in2(N__20166),
            .in3(N__20115),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__47478),
            .ce(),
            .sr(N__47088));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__21117),
            .in2(N__21108),
            .in3(N__21045),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__47478),
            .ce(),
            .sr(N__47088));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__21042),
            .in2(N__21036),
            .in3(N__20973),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__47478),
            .ce(),
            .sr(N__47088));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__20970),
            .in2(N__20964),
            .in3(N__20895),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__47478),
            .ce(),
            .sr(N__47088));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5  (
            .in0(_gnd_net_),
            .in1(N__20892),
            .in2(N__20883),
            .in3(N__20811),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__47478),
            .ce(),
            .sr(N__47088));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__20808),
            .in2(N__20802),
            .in3(N__20733),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__47478),
            .ce(),
            .sr(N__47088));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7  (
            .in0(_gnd_net_),
            .in1(N__22839),
            .in2(N__20730),
            .in3(N__20658),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__47478),
            .ce(),
            .sr(N__47088));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__23046),
            .in2(N__20655),
            .in3(N__20586),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__47466),
            .ce(),
            .sr(N__47090));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__21561),
            .in2(N__21552),
            .in3(N__21510),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__47466),
            .ce(),
            .sr(N__47090));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(N__21507),
            .in2(N__21498),
            .in3(N__21444),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__47466),
            .ce(),
            .sr(N__47090));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__21435),
            .in2(N__22134),
            .in3(N__21384),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__47466),
            .ce(),
            .sr(N__47090));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(N__21381),
            .in2(N__21372),
            .in3(N__21312),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__47466),
            .ce(),
            .sr(N__47090));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(N__21301),
            .in2(N__22193),
            .in3(N__21258),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__47466),
            .ce(),
            .sr(N__47090));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__22157),
            .in2(N__21255),
            .in3(N__21213),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__47466),
            .ce(),
            .sr(N__47090));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__21208),
            .in2(N__22194),
            .in3(N__21168),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__47466),
            .ce(),
            .sr(N__47090));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__22195),
            .in2(N__21165),
            .in3(N__21120),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__47458),
            .ce(),
            .sr(N__47093));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__21864),
            .in2(N__22224),
            .in3(N__21828),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__47458),
            .ce(),
            .sr(N__47093));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__22199),
            .in2(N__21825),
            .in3(N__21783),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__47458),
            .ce(),
            .sr(N__47093));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__22791),
            .in2(N__22225),
            .in3(N__21780),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__47458),
            .ce(),
            .sr(N__47093));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__22203),
            .in2(N__22751),
            .in3(N__21777),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__47458),
            .ce(),
            .sr(N__47093));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__21774),
            .in2(N__22226),
            .in3(N__21735),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__47458),
            .ce(),
            .sr(N__47093));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__22207),
            .in2(N__21732),
            .in3(N__21672),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__47458),
            .ce(),
            .sr(N__47093));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__22833),
            .in2(N__22227),
            .in3(N__21654),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__47458),
            .ce(),
            .sr(N__47093));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__21650),
            .in2(N__22228),
            .in3(N__21612),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__47449),
            .ce(),
            .sr(N__47094));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__22214),
            .in2(N__21609),
            .in3(N__21564),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__47449),
            .ce(),
            .sr(N__47094));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__22122),
            .in2(N__22229),
            .in3(N__22083),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__47449),
            .ce(),
            .sr(N__47094));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__22218),
            .in2(N__22080),
            .in3(N__22038),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__47449),
            .ce(),
            .sr(N__47094));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__22035),
            .in2(N__22230),
            .in3(N__21996),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__47449),
            .ce(),
            .sr(N__47094));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5  (
            .in0(_gnd_net_),
            .in1(N__22222),
            .in2(N__21993),
            .in3(N__21957),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__47449),
            .ce(),
            .sr(N__47094));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6  (
            .in0(N__22223),
            .in1(N__22707),
            .in2(_gnd_net_),
            .in3(N__21954),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47449),
            .ce(),
            .sr(N__47094));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22848),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47449),
            .ce(),
            .sr(N__47094));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_21_0  (
            .in0(N__22251),
            .in1(N__21939),
            .in2(N__22266),
            .in3(N__21924),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_21_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_21_1  (
            .in0(N__22290),
            .in1(N__21903),
            .in2(N__21891),
            .in3(N__22302),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_21_2  (
            .in0(N__22353),
            .in1(N__22403),
            .in2(N__22365),
            .in3(N__22388),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_3_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_3_21_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_3_21_3  (
            .in0(_gnd_net_),
            .in1(N__22364),
            .in2(_gnd_net_),
            .in3(N__22352),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_3_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_3_21_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_3_21_4  (
            .in0(N__22344),
            .in1(N__22325),
            .in2(N__22311),
            .in3(N__22278),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_21_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_21_6  (
            .in0(N__22301),
            .in1(N__22289),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_21_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_21_7  (
            .in0(N__22277),
            .in1(N__22262),
            .in2(N__22254),
            .in3(N__22250),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_4_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_4_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_4_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22511),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47479),
            .ce(),
            .sr(N__47081));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_4_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_4_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23091),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47479),
            .ce(),
            .sr(N__47081));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22892),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47479),
            .ce(),
            .sr(N__47081));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_4_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24380),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47467),
            .ce(),
            .sr(N__47085));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22973),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47467),
            .ce(),
            .sr(N__47085));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_18_2  (
            .in0(N__22832),
            .in1(N__22790),
            .in2(N__22752),
            .in3(N__22697),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__22545),
            .in2(_gnd_net_),
            .in3(N__24114),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_5_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_5_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__24105),
            .in2(_gnd_net_),
            .in3(N__22521),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__47480),
            .ce(),
            .sr(N__47073));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_5_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_5_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__24348),
            .in2(_gnd_net_),
            .in3(N__22497),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__47480),
            .ce(),
            .sr(N__47073));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_5_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_5_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__24336),
            .in2(_gnd_net_),
            .in3(N__22470),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__47480),
            .ce(),
            .sr(N__47073));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_5_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_5_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__24324),
            .in2(_gnd_net_),
            .in3(N__22437),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__47480),
            .ce(),
            .sr(N__47073));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_5_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_5_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_5_15_5  (
            .in0(_gnd_net_),
            .in1(N__24312),
            .in2(_gnd_net_),
            .in3(N__22407),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__47480),
            .ce(),
            .sr(N__47073));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_5_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_5_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_5_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(N__24300),
            .in2(_gnd_net_),
            .in3(N__23007),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__47480),
            .ce(),
            .sr(N__47073));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_5_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_5_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_5_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(N__24288),
            .in2(_gnd_net_),
            .in3(N__22980),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__47480),
            .ce(),
            .sr(N__47073));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_5_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_5_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_5_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(N__24276),
            .in2(_gnd_net_),
            .in3(N__22959),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_5_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__47468),
            .ce(),
            .sr(N__47076));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_5_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_5_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_5_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(N__24264),
            .in2(_gnd_net_),
            .in3(N__22956),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__47468),
            .ce(),
            .sr(N__47076));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_5_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_5_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_5_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(N__24447),
            .in2(_gnd_net_),
            .in3(N__22929),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__47468),
            .ce(),
            .sr(N__47076));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_5_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_5_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(N__24435),
            .in2(_gnd_net_),
            .in3(N__22902),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__47468),
            .ce(),
            .sr(N__47076));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_5_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_5_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_5_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(N__24423),
            .in2(_gnd_net_),
            .in3(N__22878),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__47468),
            .ce(),
            .sr(N__47076));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_5_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_5_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_5_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_5_16_5  (
            .in0(_gnd_net_),
            .in1(N__23352),
            .in2(_gnd_net_),
            .in3(N__22851),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__47468),
            .ce(),
            .sr(N__47076));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_5_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_5_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(N__24408),
            .in2(_gnd_net_),
            .in3(N__23163),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47468),
            .ce(),
            .sr(N__47076));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23066),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47450),
            .ce(),
            .sr(N__47086));
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_7_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_7_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_7_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_23_LC_7_7_5  (
            .in0(N__26514),
            .in1(N__26539),
            .in2(_gnd_net_),
            .in3(N__41184),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47548),
            .ce(N__32100),
            .sr(N__47029));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_7_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_7_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_7_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_7_8_6  (
            .in0(N__41133),
            .in1(N__24961),
            .in2(_gnd_net_),
            .in3(N__24940),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47540),
            .ce(N__32112),
            .sr(N__47035));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_7_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_7_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_7_8_7  (
            .in0(N__25093),
            .in1(N__25068),
            .in2(_gnd_net_),
            .in3(N__41132),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_7_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_7_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_7_9_5  (
            .in0(N__25015),
            .in1(N__24980),
            .in2(_gnd_net_),
            .in3(N__41181),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(elapsed_time_ns_1_RNI02CN9_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_7_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_7_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_7_9_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_7_9_6  (
            .in0(N__41182),
            .in1(_gnd_net_),
            .in2(N__23037),
            .in3(N__25016),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47531),
            .ce(N__32101),
            .sr(N__47041));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__23653),
            .in2(N__23703),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47519),
            .ce(N__25221),
            .sr(N__47046));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__23632),
            .in2(N__23679),
            .in3(N__23034),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47519),
            .ce(N__25221),
            .sr(N__47046));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__23654),
            .in2(N__23612),
            .in3(N__23193),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47519),
            .ce(N__25221),
            .sr(N__47046));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(N__23584),
            .in2(N__23637),
            .in3(N__23190),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47519),
            .ce(N__25221),
            .sr(N__47046));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__23563),
            .in2(N__23613),
            .in3(N__23187),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47519),
            .ce(N__25221),
            .sr(N__47046));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__23887),
            .in2(N__23589),
            .in3(N__23184),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47519),
            .ce(N__25221),
            .sr(N__47046));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__23564),
            .in2(N__23871),
            .in3(N__23181),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47519),
            .ce(N__25221),
            .sr(N__47046));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__23888),
            .in2(N__23841),
            .in3(N__23178),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47519),
            .ce(N__25221),
            .sr(N__47046));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__23809),
            .in2(N__23870),
            .in3(N__23175),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47506),
            .ce(N__25220),
            .sr(N__47052));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__23788),
            .in2(N__23840),
            .in3(N__23172),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47506),
            .ce(N__25220),
            .sr(N__47052));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__23810),
            .in2(N__23768),
            .in3(N__23169),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47506),
            .ce(N__25220),
            .sr(N__47052));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__23740),
            .in2(N__23793),
            .in3(N__23166),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47506),
            .ce(N__25220),
            .sr(N__47052));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__23719),
            .in2(N__23769),
            .in3(N__23220),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47506),
            .ce(N__25220),
            .sr(N__47052));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__24091),
            .in2(N__23745),
            .in3(N__23217),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47506),
            .ce(N__25220),
            .sr(N__47052));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__23720),
            .in2(N__24075),
            .in3(N__23214),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47506),
            .ce(N__25220),
            .sr(N__47052));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__24092),
            .in2(N__24045),
            .in3(N__23211),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47506),
            .ce(N__25220),
            .sr(N__47052));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__24013),
            .in2(N__24074),
            .in3(N__23208),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47493),
            .ce(N__25218),
            .sr(N__47056));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__23992),
            .in2(N__24044),
            .in3(N__23205),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47493),
            .ce(N__25218),
            .sr(N__47056));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__24014),
            .in2(N__23972),
            .in3(N__23202),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47493),
            .ce(N__25218),
            .sr(N__47056));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__23944),
            .in2(N__23997),
            .in3(N__23199),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47493),
            .ce(N__25218),
            .sr(N__47056));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__23923),
            .in2(N__23973),
            .in3(N__23196),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47493),
            .ce(N__25218),
            .sr(N__47056));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__23905),
            .in2(N__23949),
            .in3(N__23244),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47493),
            .ce(N__25218),
            .sr(N__47056));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(N__23924),
            .in2(N__24252),
            .in3(N__23241),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47493),
            .ce(N__25218),
            .sr(N__47056));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__23906),
            .in2(N__24222),
            .in3(N__23238),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47493),
            .ce(N__25218),
            .sr(N__47056));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__24187),
            .in2(N__24251),
            .in3(N__23235),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47481),
            .ce(N__25217),
            .sr(N__47059));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__24163),
            .in2(N__24221),
            .in3(N__23232),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47481),
            .ce(N__25217),
            .sr(N__47059));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__24143),
            .in2(N__24192),
            .in3(N__23229),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47481),
            .ce(N__25217),
            .sr(N__47059));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__24125),
            .in2(N__24168),
            .in3(N__23226),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47481),
            .ce(N__25217),
            .sr(N__47059));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23223),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47481),
            .ce(N__25217),
            .sr(N__47059));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_7_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_7_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_7_14_0  (
            .in0(N__25906),
            .in1(N__25867),
            .in2(_gnd_net_),
            .in3(N__41169),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_7_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_7_16_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_7_16_0  (
            .in0(N__25395),
            .in1(N__41196),
            .in2(_gnd_net_),
            .in3(N__25416),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47451),
            .ce(N__32111),
            .sr(N__47068));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_7_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_7_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24404),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42407),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_7_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_7_25_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_7_25_6  (
            .in0(N__27307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27269),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_7_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_7_26_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_7_26_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23328),
            .in3(N__23343),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_7_26_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_7_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_7_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_7_26_1  (
            .in0(_gnd_net_),
            .in1(N__23307),
            .in2(_gnd_net_),
            .in3(N__23319),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_7_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_7_26_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_7_26_2  (
            .in0(_gnd_net_),
            .in1(N__23286),
            .in2(_gnd_net_),
            .in3(N__23301),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_7_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_7_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_7_26_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_7_26_3  (
            .in0(_gnd_net_),
            .in1(N__23265),
            .in2(_gnd_net_),
            .in3(N__23280),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_7_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_7_26_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_7_26_4  (
            .in0(_gnd_net_),
            .in1(N__23469),
            .in2(_gnd_net_),
            .in3(N__23259),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_7_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_7_26_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_7_26_5  (
            .in0(_gnd_net_),
            .in1(N__23448),
            .in2(_gnd_net_),
            .in3(N__23463),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_7_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_7_26_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_7_26_6  (
            .in0(_gnd_net_),
            .in1(N__23427),
            .in2(_gnd_net_),
            .in3(N__23442),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_7_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_7_26_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_7_26_7  (
            .in0(_gnd_net_),
            .in1(N__23406),
            .in2(_gnd_net_),
            .in3(N__23421),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_7_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_7_27_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_7_27_0  (
            .in0(_gnd_net_),
            .in1(N__23385),
            .in2(_gnd_net_),
            .in3(N__23400),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_7_27_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_7_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_7_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_7_27_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_7_27_1  (
            .in0(N__23379),
            .in1(N__23367),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_7_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_7_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_7_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_7_27_2  (
            .in0(_gnd_net_),
            .in1(N__27308),
            .in2(_gnd_net_),
            .in3(N__23361),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_7_27_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_7_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_7_27_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_7_27_3  (
            .in0(N__29873),
            .in1(N__25649),
            .in2(_gnd_net_),
            .in3(N__23358),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_7_27_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_7_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_7_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_7_27_4  (
            .in0(_gnd_net_),
            .in1(N__29932),
            .in2(_gnd_net_),
            .in3(N__23355),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_7_27_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_7_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_7_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_7_27_5  (
            .in0(_gnd_net_),
            .in1(N__27226),
            .in2(_gnd_net_),
            .in3(N__23499),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_7_27_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_7_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_7_27_6  (
            .in0(_gnd_net_),
            .in1(N__27325),
            .in2(_gnd_net_),
            .in3(N__23496),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_7_27_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_7_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_7_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_7_27_7  (
            .in0(_gnd_net_),
            .in1(N__29776),
            .in2(_gnd_net_),
            .in3(N__23493),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_7_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_7_28_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_7_28_0  (
            .in0(_gnd_net_),
            .in1(N__27388),
            .in2(_gnd_net_),
            .in3(N__23490),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_7_28_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_7_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_7_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_7_28_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_7_28_1  (
            .in0(_gnd_net_),
            .in1(N__27427),
            .in2(_gnd_net_),
            .in3(N__23487),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_7_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_7_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_7_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_7_28_2  (
            .in0(_gnd_net_),
            .in1(N__25699),
            .in2(_gnd_net_),
            .in3(N__23484),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_7_28_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_7_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_7_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_7_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23481),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23478),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47552),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_8_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_8_7_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_8_7_0  (
            .in0(N__28295),
            .in1(N__23523),
            .in2(N__28323),
            .in3(N__23511),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_8_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_8_7_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_8_7_1  (
            .in0(N__23510),
            .in1(N__28322),
            .in2(N__28299),
            .in3(N__23522),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_8_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_8_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_8_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_22_LC_8_7_5  (
            .in0(N__26624),
            .in1(N__26590),
            .in2(_gnd_net_),
            .in3(N__41138),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47541),
            .ce(N__32106),
            .sr(N__47023));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_8_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_8_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_8_8_0  (
            .in0(N__26170),
            .in1(N__26217),
            .in2(N__25071),
            .in3(N__26286),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_8_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_8_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_8_8_1  (
            .in0(N__23547),
            .in1(N__23535),
            .in2(N__23502),
            .in3(N__23529),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_8_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__25384),
            .in2(_gnd_net_),
            .in3(N__26046),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_8_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_8_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_8_8_3  (
            .in0(N__24965),
            .in1(N__24939),
            .in2(_gnd_net_),
            .in3(N__41135),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_8_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_8_8_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_8_8_4  (
            .in0(N__24612),
            .in1(N__26355),
            .in2(_gnd_net_),
            .in3(N__23541),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_8_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_8_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_8_8_5  (
            .in0(N__24581),
            .in1(N__24613),
            .in2(_gnd_net_),
            .in3(N__41136),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_8_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_8_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_8_8_6  (
            .in0(N__41134),
            .in1(N__26543),
            .in2(_gnd_net_),
            .in3(N__26521),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_8_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_8_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_8_9_0  (
            .in0(N__26805),
            .in1(N__24768),
            .in2(N__27080),
            .in3(N__41235),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_8_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_8_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_8_9_2  (
            .in0(N__25126),
            .in1(N__26103),
            .in2(N__24529),
            .in3(N__24840),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_9_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_9_3  (
            .in0(N__24722),
            .in1(_gnd_net_),
            .in2(N__41187),
            .in3(N__24697),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_8_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_8_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_8_9_4  (
            .in0(N__24522),
            .in1(N__41143),
            .in2(_gnd_net_),
            .in3(N__24560),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_8_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_8_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_8_9_5  (
            .in0(N__25866),
            .in1(N__26748),
            .in2(N__26523),
            .in3(N__26580),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_8_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_8_9_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_8_9_6  (
            .in0(N__26806),
            .in1(N__41142),
            .in2(_gnd_net_),
            .in3(N__26831),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_8_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_8_9_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_8_9_7  (
            .in0(N__24873),
            .in1(N__24696),
            .in2(N__24944),
            .in3(N__25011),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_10_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_10_2  (
            .in0(N__23702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47507),
            .ce(N__25219),
            .sr(N__47042));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23678),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47507),
            .ce(N__25219),
            .sr(N__47042));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_8_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_8_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_8_10_4  (
            .in0(N__24818),
            .in1(N__24841),
            .in2(_gnd_net_),
            .in3(N__41160),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_8_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_8_10_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_8_10_5  (
            .in0(N__41159),
            .in1(N__26080),
            .in2(_gnd_net_),
            .in3(N__26104),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_8_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_8_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_8_10_6  (
            .in0(N__25163),
            .in1(N__25127),
            .in2(_gnd_net_),
            .in3(N__41161),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_11_0  (
            .in0(N__25324),
            .in1(N__23698),
            .in2(_gnd_net_),
            .in3(N__23682),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__47494),
            .ce(N__25548),
            .sr(N__47047));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_11_1  (
            .in0(N__25347),
            .in1(N__23674),
            .in2(_gnd_net_),
            .in3(N__23658),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__47494),
            .ce(N__25548),
            .sr(N__47047));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_11_2  (
            .in0(N__25325),
            .in1(N__23655),
            .in2(_gnd_net_),
            .in3(N__23640),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__47494),
            .ce(N__25548),
            .sr(N__47047));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_11_3  (
            .in0(N__25348),
            .in1(N__23633),
            .in2(_gnd_net_),
            .in3(N__23616),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__47494),
            .ce(N__25548),
            .sr(N__47047));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_11_4  (
            .in0(N__25326),
            .in1(N__23611),
            .in2(_gnd_net_),
            .in3(N__23592),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__47494),
            .ce(N__25548),
            .sr(N__47047));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_11_5  (
            .in0(N__25349),
            .in1(N__23585),
            .in2(_gnd_net_),
            .in3(N__23568),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__47494),
            .ce(N__25548),
            .sr(N__47047));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_11_6  (
            .in0(N__25327),
            .in1(N__23565),
            .in2(_gnd_net_),
            .in3(N__23550),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__47494),
            .ce(N__25548),
            .sr(N__47047));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_11_7  (
            .in0(N__25350),
            .in1(N__23889),
            .in2(_gnd_net_),
            .in3(N__23874),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__47494),
            .ce(N__25548),
            .sr(N__47047));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_12_0  (
            .in0(N__25323),
            .in1(N__23863),
            .in2(_gnd_net_),
            .in3(N__23844),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__47482),
            .ce(N__25547),
            .sr(N__47053));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_12_1  (
            .in0(N__25331),
            .in1(N__23833),
            .in2(_gnd_net_),
            .in3(N__23814),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__47482),
            .ce(N__25547),
            .sr(N__47053));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_12_2  (
            .in0(N__25320),
            .in1(N__23811),
            .in2(_gnd_net_),
            .in3(N__23796),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__47482),
            .ce(N__25547),
            .sr(N__47053));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_12_3  (
            .in0(N__25328),
            .in1(N__23789),
            .in2(_gnd_net_),
            .in3(N__23772),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__47482),
            .ce(N__25547),
            .sr(N__47053));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_12_4  (
            .in0(N__25321),
            .in1(N__23767),
            .in2(_gnd_net_),
            .in3(N__23748),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__47482),
            .ce(N__25547),
            .sr(N__47053));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_12_5  (
            .in0(N__25329),
            .in1(N__23741),
            .in2(_gnd_net_),
            .in3(N__23724),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__47482),
            .ce(N__25547),
            .sr(N__47053));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_12_6  (
            .in0(N__25322),
            .in1(N__23721),
            .in2(_gnd_net_),
            .in3(N__23706),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__47482),
            .ce(N__25547),
            .sr(N__47053));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_12_7  (
            .in0(N__25330),
            .in1(N__24093),
            .in2(_gnd_net_),
            .in3(N__24078),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__47482),
            .ce(N__25547),
            .sr(N__47053));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_13_0  (
            .in0(N__25316),
            .in1(N__24067),
            .in2(_gnd_net_),
            .in3(N__24048),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__47469),
            .ce(N__25546),
            .sr(N__47057));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_13_1  (
            .in0(N__25334),
            .in1(N__24037),
            .in2(_gnd_net_),
            .in3(N__24018),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__47469),
            .ce(N__25546),
            .sr(N__47057));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_13_2  (
            .in0(N__25317),
            .in1(N__24015),
            .in2(_gnd_net_),
            .in3(N__24000),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__47469),
            .ce(N__25546),
            .sr(N__47057));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_13_3  (
            .in0(N__25335),
            .in1(N__23993),
            .in2(_gnd_net_),
            .in3(N__23976),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__47469),
            .ce(N__25546),
            .sr(N__47057));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_13_4  (
            .in0(N__25318),
            .in1(N__23971),
            .in2(_gnd_net_),
            .in3(N__23952),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__47469),
            .ce(N__25546),
            .sr(N__47057));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_13_5  (
            .in0(N__25336),
            .in1(N__23945),
            .in2(_gnd_net_),
            .in3(N__23928),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__47469),
            .ce(N__25546),
            .sr(N__47057));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_13_6  (
            .in0(N__25319),
            .in1(N__23925),
            .in2(_gnd_net_),
            .in3(N__23910),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__47469),
            .ce(N__25546),
            .sr(N__47057));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_13_7  (
            .in0(N__25337),
            .in1(N__23907),
            .in2(_gnd_net_),
            .in3(N__23892),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__47469),
            .ce(N__25546),
            .sr(N__47057));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_14_0  (
            .in0(N__25312),
            .in1(N__24244),
            .in2(_gnd_net_),
            .in3(N__24225),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__47459),
            .ce(N__25536),
            .sr(N__47060));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_14_1  (
            .in0(N__25332),
            .in1(N__24214),
            .in2(_gnd_net_),
            .in3(N__24195),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__47459),
            .ce(N__25536),
            .sr(N__47060));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_14_2  (
            .in0(N__25313),
            .in1(N__24188),
            .in2(_gnd_net_),
            .in3(N__24171),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__47459),
            .ce(N__25536),
            .sr(N__47060));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_14_3  (
            .in0(N__25333),
            .in1(N__24164),
            .in2(_gnd_net_),
            .in3(N__24147),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__47459),
            .ce(N__25536),
            .sr(N__47060));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_14_4  (
            .in0(N__25314),
            .in1(N__24144),
            .in2(_gnd_net_),
            .in3(N__24132),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__47459),
            .ce(N__25536),
            .sr(N__47060));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_14_5  (
            .in0(N__24126),
            .in1(N__25315),
            .in2(_gnd_net_),
            .in3(N__24129),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47459),
            .ce(N__25536),
            .sr(N__47060));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_8_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_8_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__25496),
            .in2(N__25473),
            .in3(N__25471),
            .lcout(\current_shift_inst.control_input_18 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_15_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__25503),
            .in2(_gnd_net_),
            .in3(N__24096),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__25485),
            .in2(_gnd_net_),
            .in3(N__24339),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_15_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__25479),
            .in2(_gnd_net_),
            .in3(N__24327),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_15_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__29418),
            .in2(_gnd_net_),
            .in3(N__24315),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__25452),
            .in2(_gnd_net_),
            .in3(N__24303),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_15_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__29439),
            .in2(_gnd_net_),
            .in3(N__24291),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_15_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__25446),
            .in2(_gnd_net_),
            .in3(N__24279),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_16_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__26949),
            .in2(_gnd_net_),
            .in3(N__24267),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_16_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(N__26937),
            .in2(_gnd_net_),
            .in3(N__24255),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_16_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(N__26925),
            .in2(_gnd_net_),
            .in3(N__24438),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_16_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(N__29457),
            .in2(_gnd_net_),
            .in3(N__24426),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_16_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__24393),
            .in2(_gnd_net_),
            .in3(N__24414),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_8_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_8_16_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(N__35298),
            .in2(_gnd_net_),
            .in3(N__24411),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35297),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__25497),
            .in2(_gnd_net_),
            .in3(N__25472),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47437),
            .ce(),
            .sr(N__47069));
    defparam \phase_controller_inst2.S2_LC_8_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_8_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_8_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_8_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41955),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47424),
            .ce(),
            .sr(N__47091));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_8_26_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_8_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_8_26_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_8_26_2  (
            .in0(N__27329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27344),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_8_26_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_8_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_8_26_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_8_26_7  (
            .in0(N__27230),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27248),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_8_27_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_8_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_8_27_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_8_27_2  (
            .in0(N__29780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29753),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_8_27_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_8_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_8_27_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_8_27_3  (
            .in0(N__27371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27392),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_8_27_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_8_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_8_27_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_8_27_4  (
            .in0(_gnd_net_),
            .in1(N__29906),
            .in2(_gnd_net_),
            .in3(N__29936),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_8_27_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_8_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_8_27_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_8_27_5  (
            .in0(_gnd_net_),
            .in1(N__27446),
            .in2(_gnd_net_),
            .in3(N__27431),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_8_27_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_8_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_8_27_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_8_27_6  (
            .in0(N__25700),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25712),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_5.C_ON=1'b0;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47559),
            .lcout(GB_BUFFER_clock_output_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_6.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_6 (
            .in0(N__24471),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_9_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_9_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_9_4_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_25_LC_9_4_6  (
            .in0(N__27097),
            .in1(N__27079),
            .in2(_gnd_net_),
            .in3(N__41183),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47553),
            .ce(N__32071),
            .sr(N__46996));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_9_5_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_9_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_9_5_0  (
            .in0(N__24797),
            .in1(N__24776),
            .in2(_gnd_net_),
            .in3(N__41137),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_9_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_9_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_9_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_26_LC_9_6_6  (
            .in0(N__41109),
            .in1(N__24793),
            .in2(_gnd_net_),
            .in3(N__24777),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47542),
            .ce(N__32018),
            .sr(N__47010));
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_9_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_9_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_9_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_24_LC_9_6_7  (
            .in0(N__26763),
            .in1(N__26717),
            .in2(_gnd_net_),
            .in3(N__41110),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47542),
            .ce(N__32018),
            .sr(N__47010));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0  (
            .in0(N__28430),
            .in1(N__28406),
            .in2(N__24498),
            .in3(N__24486),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_7_1  (
            .in0(N__40949),
            .in1(N__24905),
            .in2(_gnd_net_),
            .in3(N__24883),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_3 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_3  (
            .in0(N__24485),
            .in1(N__28431),
            .in2(N__28410),
            .in3(N__24494),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_7_4  (
            .in0(N__26177),
            .in1(N__26138),
            .in2(_gnd_net_),
            .in3(N__40950),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(elapsed_time_ns_1_RNI68CN9_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_7_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_9_7_5  (
            .in0(N__40951),
            .in1(_gnd_net_),
            .in2(N__24501),
            .in3(N__26178),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47532),
            .ce(N__32105),
            .sr(N__47016));
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_9_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_9_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_9_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_28_LC_9_8_1  (
            .in0(N__24621),
            .in1(N__24577),
            .in2(_gnd_net_),
            .in3(N__40993),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47520),
            .ce(N__32107),
            .sr(N__47024));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_8_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_9_8_2  (
            .in0(N__40991),
            .in1(N__26239),
            .in2(_gnd_net_),
            .in3(N__26222),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47520),
            .ce(N__32107),
            .sr(N__47024));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_8_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__40992),
            .in2(N__26685),
            .in3(N__26661),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47520),
            .ce(N__32107),
            .sr(N__47024));
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_9_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_9_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_9_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_29_LC_9_8_5  (
            .in0(N__26827),
            .in1(N__26811),
            .in2(_gnd_net_),
            .in3(N__40994),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47520),
            .ce(N__32107),
            .sr(N__47024));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_9_8_6  (
            .in0(N__40990),
            .in1(N__24901),
            .in2(_gnd_net_),
            .in3(N__24885),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47520),
            .ce(N__32107),
            .sr(N__47024));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_9_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_9_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_9_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_9_8_7  (
            .in0(N__25787),
            .in1(N__25981),
            .in2(_gnd_net_),
            .in3(N__40995),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47520),
            .ce(N__32107),
            .sr(N__47024));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_9_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_9_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_9_9_0  (
            .in0(N__40996),
            .in1(N__24814),
            .in2(_gnd_net_),
            .in3(N__24842),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47508),
            .ce(N__32079),
            .sr(N__47030));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_9_9_1  (
            .in0(N__24637),
            .in1(N__24668),
            .in2(_gnd_net_),
            .in3(N__40999),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47508),
            .ce(N__32079),
            .sr(N__47030));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_9_9_2  (
            .in0(N__40998),
            .in1(N__24556),
            .in2(_gnd_net_),
            .in3(N__24540),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47508),
            .ce(N__32079),
            .sr(N__47030));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_9_9_3  (
            .in0(N__24718),
            .in1(N__24702),
            .in2(_gnd_net_),
            .in3(N__41000),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47508),
            .ce(N__32079),
            .sr(N__47030));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_9_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_9_9_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_9_9_4  (
            .in0(N__40997),
            .in1(N__25159),
            .in2(_gnd_net_),
            .in3(N__25139),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47508),
            .ce(N__32079),
            .sr(N__47030));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_7  (
            .in0(N__25100),
            .in1(N__25070),
            .in2(_gnd_net_),
            .in3(N__41001),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47508),
            .ce(N__32079),
            .sr(N__47030));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0  (
            .in0(N__26424),
            .in1(N__26390),
            .in2(N__26664),
            .in3(N__24660),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2  (
            .in0(N__24639),
            .in1(N__24661),
            .in2(_gnd_net_),
            .in3(N__41162),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6  (
            .in0(N__26425),
            .in1(N__26459),
            .in2(_gnd_net_),
            .in3(N__41163),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47495),
            .ce(N__32070),
            .sr(N__47036));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7  (
            .in0(N__26391),
            .in1(N__41167),
            .in2(_gnd_net_),
            .in3(N__26406),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47495),
            .ce(N__32070),
            .sr(N__47036));
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_9_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_9_11_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_26_LC_9_11_0  (
            .in0(N__24798),
            .in1(N__24772),
            .in2(_gnd_net_),
            .in3(N__41127),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47483),
            .ce(N__27019),
            .sr(N__47043));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_9_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_9_11_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_9_11_1  (
            .in0(N__41121),
            .in1(N__24726),
            .in2(_gnd_net_),
            .in3(N__24701),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47483),
            .ce(N__27019),
            .sr(N__47043));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_9_11_2  (
            .in0(N__24669),
            .in1(N__24638),
            .in2(_gnd_net_),
            .in3(N__41125),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47483),
            .ce(N__27019),
            .sr(N__47043));
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_9_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_9_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_28_LC_9_11_3  (
            .in0(N__41122),
            .in1(N__24620),
            .in2(_gnd_net_),
            .in3(N__24582),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47483),
            .ce(N__27019),
            .sr(N__47043));
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_9_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_9_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_21_LC_9_11_4  (
            .in0(N__25907),
            .in1(N__25874),
            .in2(_gnd_net_),
            .in3(N__41126),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47483),
            .ce(N__27019),
            .sr(N__47043));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_9_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_9_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_9_11_5  (
            .in0(N__41124),
            .in1(N__26013),
            .in2(_gnd_net_),
            .in3(N__26057),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47483),
            .ce(N__27019),
            .sr(N__47043));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_9_11_6  (
            .in0(N__24561),
            .in1(N__24536),
            .in2(_gnd_net_),
            .in3(N__41128),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47483),
            .ce(N__27019),
            .sr(N__47043));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_9_11_7  (
            .in0(N__41123),
            .in1(N__25164),
            .in2(_gnd_net_),
            .in3(N__25143),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47483),
            .ce(N__27019),
            .sr(N__47043));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_12_0 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_12_0  (
            .in0(N__31089),
            .in1(N__25110),
            .in2(N__25029),
            .in3(N__31112),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_12_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_12_1  (
            .in0(N__25109),
            .in1(N__31088),
            .in2(N__31116),
            .in3(N__25025),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_9_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_9_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_9_12_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_9_12_3  (
            .in0(N__25101),
            .in1(N__41179),
            .in2(_gnd_net_),
            .in3(N__25069),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47470),
            .ce(N__27017),
            .sr(N__47048));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_9_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_9_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_9_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_9_12_4  (
            .in0(N__25017),
            .in1(N__24987),
            .in2(_gnd_net_),
            .in3(N__41165),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47470),
            .ce(N__27017),
            .sr(N__47048));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_9_12_5  (
            .in0(N__41164),
            .in1(N__24969),
            .in2(_gnd_net_),
            .in3(N__24945),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47470),
            .ce(N__27017),
            .sr(N__47048));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_9_12_6  (
            .in0(N__24906),
            .in1(N__24884),
            .in2(_gnd_net_),
            .in3(N__41166),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47470),
            .ce(N__27017),
            .sr(N__47048));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_9_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_9_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_9_12_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_9_12_7  (
            .in0(N__24846),
            .in1(N__41180),
            .in2(_gnd_net_),
            .in3(N__24819),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47470),
            .ce(N__27017),
            .sr(N__47048));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_13_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_13_0  (
            .in0(N__31016),
            .in1(N__30989),
            .in2(N__25440),
            .in3(N__25425),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_13_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_13_1  (
            .in0(N__25424),
            .in1(N__31017),
            .in2(N__30993),
            .in3(N__25436),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_9_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_9_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_9_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_20_LC_9_13_2  (
            .in0(N__41190),
            .in1(N__26289),
            .in2(_gnd_net_),
            .in3(N__25833),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47460),
            .ce(N__27015),
            .sr(N__47054));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_9_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_9_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_9_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_9_13_4  (
            .in0(N__41191),
            .in1(N__25982),
            .in2(_gnd_net_),
            .in3(N__25794),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47460),
            .ce(N__27015),
            .sr(N__47054));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_5  (
            .in0(N__25393),
            .in1(N__41189),
            .in2(_gnd_net_),
            .in3(N__25409),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(elapsed_time_ns_1_RNIK63T9_0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_9_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_9_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_9_13_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_9_13_6  (
            .in0(N__41192),
            .in1(_gnd_net_),
            .in2(N__25398),
            .in3(N__25394),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47460),
            .ce(N__27015),
            .sr(N__47054));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_14_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_14_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_9_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25362),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47452),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_9_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_9_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_9_14_3  (
            .in0(N__41170),
            .in1(N__26356),
            .in2(_gnd_net_),
            .in3(N__26311),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_9_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_9_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26964),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_14_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_14_5  (
            .in0(N__26966),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28142),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_198_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_14_6 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__26965),
            .in2(N__28146),
            .in3(N__29732),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_199_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_15_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_15_0  (
            .in0(N__26458),
            .in1(N__26436),
            .in2(_gnd_net_),
            .in3(N__41188),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_16_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_16_0  (
            .in0(N__35286),
            .in1(N__31578),
            .in2(_gnd_net_),
            .in3(N__29367),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_9_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_9_16_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_9_16_1  (
            .in0(N__31593),
            .in1(N__29256),
            .in2(_gnd_net_),
            .in3(N__35284),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_9_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_9_16_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_9_16_2  (
            .in0(N__35287),
            .in1(N__31563),
            .in2(_gnd_net_),
            .in3(N__29352),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_16_3 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_16_3  (
            .in0(N__31548),
            .in1(N__29337),
            .in2(_gnd_net_),
            .in3(N__35288),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_16_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_16_4  (
            .in0(N__35285),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.N_1288_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_9_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_9_16_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_9_16_5  (
            .in0(N__31680),
            .in1(N__29319),
            .in2(_gnd_net_),
            .in3(N__35289),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_9_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_9_16_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_9_16_7  (
            .in0(N__31653),
            .in1(N__29301),
            .in2(_gnd_net_),
            .in3(N__35290),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0  (
            .in0(_gnd_net_),
            .in1(N__25650),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_26_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1  (
            .in0(_gnd_net_),
            .in1(N__25617),
            .in2(_gnd_net_),
            .in3(N__25602),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2  (
            .in0(_gnd_net_),
            .in1(N__25599),
            .in2(_gnd_net_),
            .in3(N__25584),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3  (
            .in0(_gnd_net_),
            .in1(N__25581),
            .in2(_gnd_net_),
            .in3(N__25566),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4  (
            .in0(_gnd_net_),
            .in1(N__27159),
            .in2(_gnd_net_),
            .in3(N__25563),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5  (
            .in0(_gnd_net_),
            .in1(N__35467),
            .in2(N__27114),
            .in3(N__25560),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6  (
            .in0(_gnd_net_),
            .in1(N__27798),
            .in2(N__35538),
            .in3(N__25557),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7  (
            .in0(_gnd_net_),
            .in1(N__35471),
            .in2(N__27753),
            .in3(N__25554),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__27699),
            .in2(_gnd_net_),
            .in3(N__25551),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1  (
            .in0(_gnd_net_),
            .in1(N__27651),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2  (
            .in0(_gnd_net_),
            .in1(N__27606),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(N__27567),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4  (
            .in0(_gnd_net_),
            .in1(N__27522),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(N__28071),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6  (
            .in0(_gnd_net_),
            .in1(N__28041),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7  (
            .in0(_gnd_net_),
            .in1(N__28014),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(N__27984),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_28_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1  (
            .in0(_gnd_net_),
            .in1(N__27954),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(N__27924),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3  (
            .in0(_gnd_net_),
            .in1(N__27858),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25719),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_9_28_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_9_28_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_9_28_6 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_9_28_6  (
            .in0(N__25716),
            .in1(N__29831),
            .in2(N__25701),
            .in3(N__25680),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_5_0 .LUT_INIT=16'b0111001100010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_5_0  (
            .in0(N__28272),
            .in1(N__28250),
            .in2(N__25662),
            .in3(N__25671),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1 .LUT_INIT=16'b1000111010101111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1  (
            .in0(N__25670),
            .in1(N__25658),
            .in2(N__28251),
            .in3(N__28271),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_10_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_10_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_10_5_2  (
            .in0(N__27101),
            .in1(N__27081),
            .in2(_gnd_net_),
            .in3(N__41092),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5  (
            .in0(N__41093),
            .in1(N__29681),
            .in2(_gnd_net_),
            .in3(N__29635),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_6_0 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_6_0  (
            .in0(N__25812),
            .in1(N__28226),
            .in2(N__28562),
            .in3(N__25803),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_10_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_10_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_27_LC_10_6_3  (
            .in0(N__26364),
            .in1(N__26319),
            .in2(_gnd_net_),
            .in3(N__41105),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47521),
            .ce(N__32049),
            .sr(N__46997));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_6_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_6_4  (
            .in0(N__25811),
            .in1(N__28227),
            .in2(N__28563),
            .in3(N__25802),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_6_5  (
            .in0(N__25786),
            .in1(N__25983),
            .in2(_gnd_net_),
            .in3(N__41104),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_7_0 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_7_0  (
            .in0(N__25755),
            .in1(N__28531),
            .in2(N__25767),
            .in3(N__28513),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_10_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_10_7_1 .LUT_INIT=16'b1100111101001101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_10_7_1  (
            .in0(N__28532),
            .in1(N__25766),
            .in2(N__28515),
            .in3(N__25754),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_4  (
            .in0(N__26008),
            .in1(N__26058),
            .in2(_gnd_net_),
            .in3(N__41002),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47510),
            .ce(N__32080),
            .sr(N__47005));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_8_0  (
            .in0(N__26623),
            .in1(N__26595),
            .in2(_gnd_net_),
            .in3(N__40946),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_10_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_10_8_1 .LUT_INIT=16'b1111001101110001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_10_8_1  (
            .in0(N__28187),
            .in1(N__28165),
            .in2(N__25746),
            .in3(N__25730),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_8_2 .LUT_INIT=16'b0000101010001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_8_2  (
            .in0(N__25745),
            .in1(N__25731),
            .in2(N__28167),
            .in3(N__28188),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_10_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_10_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_10_8_3  (
            .in0(N__40947),
            .in1(N__26243),
            .in2(_gnd_net_),
            .in3(N__26218),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_10_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_10_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_10_8_4  (
            .in0(N__26012),
            .in1(N__26056),
            .in2(_gnd_net_),
            .in3(N__40948),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_10_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_10_8_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_10_8_5  (
            .in0(N__25992),
            .in1(N__25977),
            .in2(N__29680),
            .in3(N__25944),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_6 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_6  (
            .in0(N__28477),
            .in1(N__25935),
            .in2(N__25926),
            .in3(N__25923),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_10_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_10_8_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(N__26758),
            .in2(N__25914),
            .in3(N__26716),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_10_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_10_9_0 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_10_9_0  (
            .in0(N__26253),
            .in1(N__25841),
            .in2(N__28385),
            .in3(N__28352),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_10_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_10_9_1 .LUT_INIT=16'b1000101011101111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_10_9_1  (
            .in0(N__25842),
            .in1(N__26252),
            .in2(N__28386),
            .in3(N__28353),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_10_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_10_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_21_LC_10_9_3  (
            .in0(N__40957),
            .in1(N__25911),
            .in2(_gnd_net_),
            .in3(N__25878),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47484),
            .ce(N__32078),
            .sr(N__47017));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_9_4  (
            .in0(N__26287),
            .in1(N__40955),
            .in2(_gnd_net_),
            .in3(N__25826),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_10_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_10_9_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_20_LC_10_9_5  (
            .in0(N__40956),
            .in1(_gnd_net_),
            .in2(N__25815),
            .in3(N__26288),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47484),
            .ce(N__32078),
            .sr(N__47017));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_10_9_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_10_9_7  (
            .in0(N__26115),
            .in1(_gnd_net_),
            .in2(N__41111),
            .in3(N__26085),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47484),
            .ce(N__32078),
            .sr(N__47017));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_10_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_10_0  (
            .in0(N__31067),
            .in1(N__31040),
            .in2(N__26127),
            .in3(N__26187),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_10_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_10_10_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_10_10_1  (
            .in0(N__26186),
            .in1(N__31068),
            .in2(N__31044),
            .in3(N__26123),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_10_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_10_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_10_10_2  (
            .in0(N__26244),
            .in1(N__26223),
            .in2(_gnd_net_),
            .in3(N__41119),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47471),
            .ce(N__27021),
            .sr(N__47025));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_10_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_10_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_10_10_3  (
            .in0(N__41115),
            .in1(N__26176),
            .in2(_gnd_net_),
            .in3(N__26142),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47471),
            .ce(N__27021),
            .sr(N__47025));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_10_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_10_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_10_10_4  (
            .in0(N__26114),
            .in1(N__26081),
            .in2(_gnd_net_),
            .in3(N__41120),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47471),
            .ce(N__27021),
            .sr(N__47025));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_10_10_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__29676),
            .in2(N__41185),
            .in3(N__29637),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47471),
            .ce(N__27021),
            .sr(N__47025));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_11_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_11_0  (
            .in0(N__31347),
            .in1(N__31370),
            .in2(N__26475),
            .in3(N__26556),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_10_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_10_11_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_10_11_1  (
            .in0(N__26555),
            .in1(N__31346),
            .in2(N__31374),
            .in3(N__26471),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_10_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_10_11_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_22_LC_10_11_2  (
            .in0(N__41096),
            .in1(N__26625),
            .in2(_gnd_net_),
            .in3(N__26594),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47461),
            .ce(N__27020),
            .sr(N__47031));
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_10_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_10_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_10_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_23_LC_10_11_3  (
            .in0(N__26547),
            .in1(N__26522),
            .in2(_gnd_net_),
            .in3(N__41098),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47461),
            .ce(N__27020),
            .sr(N__47031));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_10_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_10_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_10_11_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_10_11_4  (
            .in0(N__41097),
            .in1(N__26463),
            .in2(_gnd_net_),
            .in3(N__26435),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47461),
            .ce(N__27020),
            .sr(N__47031));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_10_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_10_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_10_11_5  (
            .in0(N__26388),
            .in1(N__26405),
            .in2(_gnd_net_),
            .in3(N__41094),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(elapsed_time_ns_1_RNIUVBN9_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_10_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_10_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_10_11_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_10_11_6  (
            .in0(N__41095),
            .in1(_gnd_net_),
            .in2(N__26394),
            .in3(N__26389),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47461),
            .ce(N__27020),
            .sr(N__47031));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_12_0 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_12_0  (
            .in0(N__26993),
            .in1(N__26979),
            .in2(N__31245),
            .in3(N__31275),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_10_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_10_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_27_LC_10_12_1  (
            .in0(N__41175),
            .in1(N__26363),
            .in2(_gnd_net_),
            .in3(N__26312),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(N__27018),
            .sr(N__47037));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_12_3 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_12_3  (
            .in0(N__26843),
            .in1(N__31184),
            .in2(N__31212),
            .in3(N__26771),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_12_4 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_12_4  (
            .in0(N__31185),
            .in1(N__31208),
            .in2(N__26775),
            .in3(N__26844),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_10_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_10_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_10_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_29_LC_10_12_5  (
            .in0(N__41176),
            .in1(N__26835),
            .in2(_gnd_net_),
            .in3(N__26807),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(N__27018),
            .sr(N__47037));
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_10_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_10_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_31_LC_10_12_6  (
            .in0(N__28488),
            .in1(N__28452),
            .in2(_gnd_net_),
            .in3(N__41178),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(N__27018),
            .sr(N__47037));
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_30_LC_10_12_7  (
            .in0(N__41177),
            .in1(N__40755),
            .in2(_gnd_net_),
            .in3(N__41242),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(N__27018),
            .sr(N__47037));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_13_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_13_0  (
            .in0(N__31296),
            .in1(N__31319),
            .in2(N__27033),
            .in3(N__26694),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_13_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_13_1  (
            .in0(N__26693),
            .in1(N__31295),
            .in2(N__31323),
            .in3(N__27029),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_10_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_10_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_10_13_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_24_LC_10_13_2  (
            .in0(N__26762),
            .in1(N__26718),
            .in2(_gnd_net_),
            .in3(N__41174),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47444),
            .ce(N__27016),
            .sr(N__47044));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_10_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_10_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_10_13_3  (
            .in0(N__41171),
            .in1(N__26662),
            .in2(_gnd_net_),
            .in3(N__26678),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(elapsed_time_ns_1_RNIV0CN9_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_10_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_10_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_10_13_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_10_13_4  (
            .in0(N__26663),
            .in1(_gnd_net_),
            .in2(N__26628),
            .in3(N__41173),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47444),
            .ce(N__27016),
            .sr(N__47044));
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_10_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_10_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_10_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_25_LC_10_13_5  (
            .in0(N__41172),
            .in1(N__27102),
            .in2(_gnd_net_),
            .in3(N__27078),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47444),
            .ce(N__27016),
            .sr(N__47044));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_13_7 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_13_7  (
            .in0(N__26994),
            .in1(N__31241),
            .in2(N__31274),
            .in3(N__26978),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_14_6 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_10_14_6  (
            .in0(N__26967),
            .in1(N__28141),
            .in2(_gnd_net_),
            .in3(N__29733),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47439),
            .ce(),
            .sr(N__47049));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_18_7  (
            .in0(N__40605),
            .in1(N__42755),
            .in2(N__40129),
            .in3(N__37134),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_10_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_10_20_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_10_20_0  (
            .in0(N__31638),
            .in1(N__29286),
            .in2(_gnd_net_),
            .in3(N__35276),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_1  (
            .in0(N__35277),
            .in1(N__31626),
            .in2(_gnd_net_),
            .in3(N__29478),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_4  (
            .in0(N__31614),
            .in1(N__29469),
            .in2(_gnd_net_),
            .in3(N__35278),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_10_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_10_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_10_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26913),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47420),
            .ce(),
            .sr(N__47082));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_2  (
            .in0(N__27915),
            .in1(N__27494),
            .in2(_gnd_net_),
            .in3(N__35884),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_3 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_3  (
            .in0(N__27495),
            .in1(N__27477),
            .in2(N__35902),
            .in3(N__27914),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_10_25_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_10_25_0 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_10_25_0  (
            .in0(N__27459),
            .in1(N__27447),
            .in2(N__29881),
            .in3(N__27435),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_10_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_10_25_2 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_10_25_2  (
            .in0(N__29868),
            .in1(N__27411),
            .in2(N__27399),
            .in3(N__27372),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_10_25_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_10_25_4 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_10_25_4  (
            .in0(N__29867),
            .in1(N__27360),
            .in2(N__27348),
            .in3(N__27333),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_10_25_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_10_25_5 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_10_25_5  (
            .in0(N__27309),
            .in1(N__27285),
            .in2(N__29880),
            .in3(N__27273),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_10_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_10_25_6 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_10_25_6  (
            .in0(N__29866),
            .in1(N__27249),
            .in2(N__27237),
            .in3(N__27210),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0  (
            .in0(_gnd_net_),
            .in1(N__27198),
            .in2(N__27180),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_10_26_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1  (
            .in0(_gnd_net_),
            .in1(N__27153),
            .in2(N__27135),
            .in3(N__27105),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2  (
            .in0(_gnd_net_),
            .in1(N__27831),
            .in2(N__27813),
            .in3(N__27792),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3  (
            .in0(_gnd_net_),
            .in1(N__27789),
            .in2(N__27774),
            .in3(N__27741),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4  (
            .in0(_gnd_net_),
            .in1(N__27738),
            .in2(N__27720),
            .in3(N__27693),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5  (
            .in0(_gnd_net_),
            .in1(N__27690),
            .in2(N__27672),
            .in3(N__27645),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6  (
            .in0(_gnd_net_),
            .in1(N__27642),
            .in2(N__27624),
            .in3(N__27600),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7  (
            .in0(_gnd_net_),
            .in1(N__27597),
            .in2(N__27585),
            .in3(N__27561),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0  (
            .in0(_gnd_net_),
            .in1(N__27558),
            .in2(N__27543),
            .in3(N__27516),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(bfn_10_27_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1  (
            .in0(_gnd_net_),
            .in1(N__27513),
            .in2(N__28095),
            .in3(N__28065),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2  (
            .in0(_gnd_net_),
            .in1(N__27908),
            .in2(N__28062),
            .in3(N__28035),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3  (
            .in0(_gnd_net_),
            .in1(N__27911),
            .in2(N__28032),
            .in3(N__28008),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4  (
            .in0(_gnd_net_),
            .in1(N__27909),
            .in2(N__28005),
            .in3(N__27978),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5  (
            .in0(_gnd_net_),
            .in1(N__27912),
            .in2(N__27975),
            .in3(N__27948),
            .lcout(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6  (
            .in0(_gnd_net_),
            .in1(N__27910),
            .in2(N__27945),
            .in3(N__27918),
            .lcout(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7  (
            .in0(_gnd_net_),
            .in1(N__27913),
            .in2(N__27870),
            .in3(N__27852),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0  (
            .in0(N__27849),
            .in1(N__27843),
            .in2(_gnd_net_),
            .in3(N__27834),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_4_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_4_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_11_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29714),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29693),
            .ce(),
            .sr(N__46975));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_5_0  (
            .in0(_gnd_net_),
            .in1(N__31830),
            .in2(N__29598),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_5_1  (
            .in0(N__32025),
            .in1(N__30071),
            .in2(_gnd_net_),
            .in3(N__28116),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__47522),
            .ce(),
            .sr(N__46981));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_5_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_5_2  (
            .in0(N__32082),
            .in1(N__30159),
            .in2(N__30035),
            .in3(N__28113),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__47522),
            .ce(),
            .sr(N__46981));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_5_3  (
            .in0(N__32026),
            .in1(N__29993),
            .in2(_gnd_net_),
            .in3(N__28110),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__47522),
            .ce(),
            .sr(N__46981));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_5_4  (
            .in0(N__32083),
            .in1(N__29969),
            .in2(_gnd_net_),
            .in3(N__28107),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__47522),
            .ce(),
            .sr(N__46981));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_5_5  (
            .in0(N__32027),
            .in1(N__30428),
            .in2(_gnd_net_),
            .in3(N__28104),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__47522),
            .ce(),
            .sr(N__46981));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_5_6  (
            .in0(N__32084),
            .in1(N__30380),
            .in2(_gnd_net_),
            .in3(N__28101),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__47522),
            .ce(),
            .sr(N__46981));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_5_7  (
            .in0(N__32028),
            .in1(N__30356),
            .in2(_gnd_net_),
            .in3(N__28098),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__47522),
            .ce(),
            .sr(N__46981));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_6_0  (
            .in0(N__32017),
            .in1(N__30296),
            .in2(_gnd_net_),
            .in3(N__28209),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__47511),
            .ce(),
            .sr(N__46989));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_6_1  (
            .in0(N__31956),
            .in1(N__30260),
            .in2(_gnd_net_),
            .in3(N__28206),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__47511),
            .ce(),
            .sr(N__46989));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_6_2  (
            .in0(N__32014),
            .in1(N__30221),
            .in2(_gnd_net_),
            .in3(N__28203),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__47511),
            .ce(),
            .sr(N__46989));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_11_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_11_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_11_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_11_6_3  (
            .in0(N__31957),
            .in1(N__30185),
            .in2(_gnd_net_),
            .in3(N__28200),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__47511),
            .ce(),
            .sr(N__46989));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_6_4  (
            .in0(N__32015),
            .in1(N__30665),
            .in2(_gnd_net_),
            .in3(N__28197),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__47511),
            .ce(),
            .sr(N__46989));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_6_5  (
            .in0(N__31958),
            .in1(N__30620),
            .in2(_gnd_net_),
            .in3(N__28194),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__47511),
            .ce(),
            .sr(N__46989));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_6_6  (
            .in0(N__32016),
            .in1(N__30578),
            .in2(_gnd_net_),
            .in3(N__28191),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__47511),
            .ce(),
            .sr(N__46989));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_6_7  (
            .in0(N__31959),
            .in1(N__28186),
            .in2(_gnd_net_),
            .in3(N__28170),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__47511),
            .ce(),
            .sr(N__46989));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_7_0  (
            .in0(N__31960),
            .in1(N__28166),
            .in2(_gnd_net_),
            .in3(N__28149),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__47497),
            .ce(),
            .sr(N__46998));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_7_1  (
            .in0(N__31964),
            .in1(N__28429),
            .in2(_gnd_net_),
            .in3(N__28413),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__47497),
            .ce(),
            .sr(N__46998));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_7_2  (
            .in0(N__31961),
            .in1(N__28405),
            .in2(_gnd_net_),
            .in3(N__28389),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__47497),
            .ce(),
            .sr(N__46998));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_11_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_11_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_11_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_11_7_3  (
            .in0(N__31965),
            .in1(N__28372),
            .in2(_gnd_net_),
            .in3(N__28356),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__47497),
            .ce(),
            .sr(N__46998));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_11_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_11_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_11_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_11_7_4  (
            .in0(N__31962),
            .in1(N__28348),
            .in2(_gnd_net_),
            .in3(N__28326),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__47497),
            .ce(),
            .sr(N__46998));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_11_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_11_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_11_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_11_7_5  (
            .in0(N__31966),
            .in1(N__28318),
            .in2(_gnd_net_),
            .in3(N__28302),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__47497),
            .ce(),
            .sr(N__46998));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_11_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_11_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_11_7_6  (
            .in0(N__31963),
            .in1(N__28294),
            .in2(_gnd_net_),
            .in3(N__28275),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__47497),
            .ce(),
            .sr(N__46998));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_11_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_11_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_11_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_11_7_7  (
            .in0(N__31967),
            .in1(N__28270),
            .in2(_gnd_net_),
            .in3(N__28254),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__47497),
            .ce(),
            .sr(N__46998));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_11_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_11_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_11_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_11_8_0  (
            .in0(N__32050),
            .in1(N__28246),
            .in2(_gnd_net_),
            .in3(N__28230),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__47485),
            .ce(),
            .sr(N__47006));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_11_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_11_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_11_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_11_8_1  (
            .in0(N__32067),
            .in1(N__28225),
            .in2(_gnd_net_),
            .in3(N__28566),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__47485),
            .ce(),
            .sr(N__47006));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_11_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_11_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_11_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_11_8_2  (
            .in0(N__32051),
            .in1(N__28555),
            .in2(_gnd_net_),
            .in3(N__28536),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__47485),
            .ce(),
            .sr(N__47006));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_11_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_11_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_11_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_11_8_3  (
            .in0(N__32068),
            .in1(N__28533),
            .in2(_gnd_net_),
            .in3(N__28518),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__47485),
            .ce(),
            .sr(N__47006));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_11_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_11_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_11_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_11_8_4  (
            .in0(N__32052),
            .in1(N__28514),
            .in2(_gnd_net_),
            .in3(N__28497),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__47485),
            .ce(),
            .sr(N__47006));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_11_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_11_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_11_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_11_8_5  (
            .in0(N__32069),
            .in1(N__28677),
            .in2(_gnd_net_),
            .in3(N__28494),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__47485),
            .ce(),
            .sr(N__47006));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_11_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_11_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_11_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_11_8_6  (
            .in0(N__32053),
            .in1(N__28646),
            .in2(_gnd_net_),
            .in3(N__28491),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47485),
            .ce(),
            .sr(N__47006));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_11_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_11_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_11_9_0  (
            .in0(N__28486),
            .in1(N__28445),
            .in2(_gnd_net_),
            .in3(N__40952),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_9_1 .LUT_INIT=16'b0100010011010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_9_1  (
            .in0(N__28658),
            .in1(N__28641),
            .in2(N__28625),
            .in3(N__28674),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_11_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_11_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_31_LC_11_9_2  (
            .in0(N__28487),
            .in1(N__28444),
            .in2(_gnd_net_),
            .in3(N__40954),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47472),
            .ce(N__32081),
            .sr(N__47011));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_9_3 .LUT_INIT=16'b1101010011011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_9_3  (
            .in0(N__28659),
            .in1(N__28645),
            .in2(N__28626),
            .in3(N__28676),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_11_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_11_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_30_LC_11_9_5  (
            .in0(N__40953),
            .in1(N__40751),
            .in2(_gnd_net_),
            .in3(N__41243),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47472),
            .ce(N__32081),
            .sr(N__47011));
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_9_6 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_9_6  (
            .in0(N__28675),
            .in1(N__28657),
            .in2(N__28647),
            .in3(N__28621),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_9_7 .LUT_INIT=16'b1111110101011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_9_7  (
            .in0(N__30136),
            .in1(N__30782),
            .in2(N__28608),
            .in3(N__30771),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_10_0 .LUT_INIT=16'b1101000011111101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_10_0  (
            .in0(N__31494),
            .in1(N__28605),
            .in2(N__31467),
            .in3(N__28589),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__32275),
            .in2(_gnd_net_),
            .in3(N__28799),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_10_2 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_10_2  (
            .in0(N__31492),
            .in1(N__28603),
            .in2(N__31466),
            .in3(N__28585),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_10_3 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_10_3  (
            .in0(N__28604),
            .in1(N__31462),
            .in2(N__28590),
            .in3(N__31493),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_hc.un4_running_df30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_10_4 .LUT_INIT=16'b1111110101011101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_10_4  (
            .in0(N__32228),
            .in1(N__29162),
            .in2(N__28572),
            .in3(N__29151),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_10_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28569),
            .in3(N__32274),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_10_6 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_10_6  (
            .in0(N__32276),
            .in1(N__32470),
            .in2(N__28803),
            .in3(N__30740),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47462),
            .ce(),
            .sr(N__47018));
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_10_7 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_11_10_7  (
            .in0(N__32229),
            .in1(N__32249),
            .in2(N__32315),
            .in3(N__32277),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47462),
            .ce(),
            .sr(N__47018));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_11_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_11_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__28791),
            .in2(N__28779),
            .in3(N__30736),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_11_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_11_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__28770),
            .in2(N__28764),
            .in3(N__30719),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_11_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_11_11_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_11_11_2  (
            .in0(N__30695),
            .in1(N__28755),
            .in2(N__28746),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_11_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_11_11_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_11_11_3  (
            .in0(N__30680),
            .in1(N__28734),
            .in2(N__28725),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_11_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_11_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__28716),
            .in2(N__28710),
            .in3(N__30965),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_11_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_11_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__28698),
            .in2(N__28686),
            .in3(N__30950),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_11_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_11_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_11_11_6  (
            .in0(N__30935),
            .in1(N__28947),
            .in2(N__28938),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_11_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_11_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__28929),
            .in2(N__28917),
            .in3(N__30920),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_11_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_11_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__28908),
            .in2(N__28902),
            .in3(N__30905),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_11_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_11_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__28893),
            .in2(N__28881),
            .in3(N__30890),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_11_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_11_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__28872),
            .in2(N__28866),
            .in3(N__30875),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_11_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_11_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__28857),
            .in2(N__28851),
            .in3(N__30860),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_11_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_11_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__28830),
            .in2(N__28842),
            .in3(N__31160),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_11_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_11_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__28821),
            .in2(N__28812),
            .in3(N__31145),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_11_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_11_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_11_12_6  (
            .in0(N__31130),
            .in1(N__29100),
            .in2(N__29112),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_11_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_11_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__29094),
            .in2(N__29082),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_11_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__29067),
            .in2(N__29055),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_11_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_11_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__29040),
            .in2(N__29031),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_11_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_11_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__29019),
            .in2(N__29010),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_11_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_11_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__28995),
            .in2(N__28989),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_11_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_11_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__28977),
            .in2(N__28971),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_11_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_11_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__28962),
            .in2(N__28956),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__29181),
            .in2(N__29169),
            .in3(N__29142),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29139),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_11_14_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_11_14_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_11_14_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_11_14_1 (
            .in0(N__29136),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47434),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__31755),
            .in2(_gnd_net_),
            .in3(N__31432),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_14_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_14_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_11_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29121),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47434),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_11_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_11_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_11_15_6 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \phase_controller_inst1.state_0_LC_11_15_6  (
            .in0(N__29202),
            .in1(N__33151),
            .in2(N__33468),
            .in3(N__32699),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47430),
            .ce(),
            .sr(N__47050));
    defparam \phase_controller_inst1.state_3_LC_11_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_11_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_11_15_7 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst1.state_3_LC_11_15_7  (
            .in0(N__31760),
            .in1(N__46388),
            .in2(N__31437),
            .in3(N__35786),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47430),
            .ce(),
            .sr(N__47050));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_11_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_11_16_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_11_16_0  (
            .in0(N__40128),
            .in1(N__40585),
            .in2(N__42852),
            .in3(N__37164),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_11_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_11_16_1 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_11_16_1  (
            .in0(N__43139),
            .in1(N__40126),
            .in2(N__40626),
            .in3(N__37379),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_11_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_11_16_2 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_11_16_2  (
            .in0(N__40125),
            .in1(N__37067),
            .in2(N__42672),
            .in3(N__40587),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_16_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_16_3  (
            .in0(N__40583),
            .in1(N__40121),
            .in2(N__46275),
            .in3(N__36885),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_11_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_11_16_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_11_16_4  (
            .in0(N__46373),
            .in1(N__40586),
            .in2(N__40229),
            .in3(N__37430),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_11_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_11_16_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_11_16_5  (
            .in0(N__40584),
            .in1(N__40127),
            .in2(N__42408),
            .in3(N__37547),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__32700),
            .in2(_gnd_net_),
            .in3(N__29201),
            .lcout(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_11_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_11_16_7 .LUT_INIT=16'b1100010111000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_11_16_7  (
            .in0(N__43281),
            .in1(N__38315),
            .in2(N__40627),
            .in3(N__40120),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__32925),
            .in2(N__33057),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__32797),
            .in2(N__31386),
            .in3(N__39444),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_17_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_17_2  (
            .in0(N__39445),
            .in1(N__39785),
            .in2(N__29190),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__39800),
            .in2(N__31416),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__39786),
            .in2(N__31395),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__39801),
            .in2(N__29241),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__39787),
            .in2(N__31512),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__39802),
            .in2(N__29229),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__39819),
            .in2(N__34632),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__29217),
            .in2(N__39972),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__39823),
            .in2(N__34728),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__29211),
            .in2(N__39973),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__39827),
            .in2(N__29277),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__31404),
            .in2(N__39974),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__39831),
            .in2(N__34602),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__29265),
            .in2(N__39975),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__39976),
            .in2(N__34713),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__34839),
            .in2(N__40133),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__39980),
            .in2(N__34686),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__34827),
            .in2(N__40134),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__39984),
            .in2(N__37287),
            .in3(N__29244),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__34815),
            .in2(N__40135),
            .in3(N__29355),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__39988),
            .in2(N__39345),
            .in3(N__29340),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__34698),
            .in2(N__40136),
            .in3(N__29325),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__40008),
            .in2(N__34659),
            .in3(N__29322),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__34803),
            .in2(N__40141),
            .in3(N__29307),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__40012),
            .in2(N__37395),
            .in3(N__29304),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__32943),
            .in2(N__40142),
            .in3(N__29289),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(N__40016),
            .in2(N__34776),
            .in3(N__29280),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(N__29487),
            .in2(N__40143),
            .in3(N__29472),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__40020),
            .in2(N__39387),
            .in3(N__29463),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_20_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_20_7  (
            .in0(N__32964),
            .in1(N__31599),
            .in2(N__35296),
            .in3(N__29460),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_11_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_11_21_2 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_11_21_2  (
            .in0(N__35283),
            .in1(_gnd_net_),
            .in2(N__31665),
            .in3(N__29445),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_11_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_11_21_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_11_21_5  (
            .in0(N__31533),
            .in1(N__29424),
            .in2(_gnd_net_),
            .in3(N__35282),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_22_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_22_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_22_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_11_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_11_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_11_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39603),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47417),
            .ce(),
            .sr(N__47077));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_11_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_11_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_11_24_0  (
            .in0(_gnd_net_),
            .in1(N__29388),
            .in2(N__29886),
            .in3(N__29885),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ),
            .ltout(),
            .carryin(bfn_11_24_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_11_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_11_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_11_24_1  (
            .in0(_gnd_net_),
            .in1(N__29382),
            .in2(_gnd_net_),
            .in3(N__29370),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_11_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_11_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(N__29895),
            .in2(_gnd_net_),
            .in3(N__29580),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_11_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_11_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(N__29577),
            .in2(_gnd_net_),
            .in3(N__29571),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_11_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_11_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_11_24_4  (
            .in0(_gnd_net_),
            .in1(N__29568),
            .in2(_gnd_net_),
            .in3(N__29562),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_11_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_11_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__29742),
            .in2(_gnd_net_),
            .in3(N__29559),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_11_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_11_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(N__29556),
            .in2(_gnd_net_),
            .in3(N__29550),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_11_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_11_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(N__29547),
            .in2(_gnd_net_),
            .in3(N__29541),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_11_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_11_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(N__29538),
            .in2(_gnd_net_),
            .in3(N__29526),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ),
            .ltout(),
            .carryin(bfn_11_25_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_11_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_11_25_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_11_25_1  (
            .in0(N__29523),
            .in1(N__29511),
            .in2(N__29872),
            .in3(N__29499),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_11_27_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_11_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_11_27_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_11_27_4  (
            .in0(N__29496),
            .in1(N__29937),
            .in2(N__29916),
            .in3(N__29829),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_11_27_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_11_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_11_27_7 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_11_27_7  (
            .in0(N__29830),
            .in1(N__29793),
            .in2(N__29784),
            .in3(N__29760),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_12_4_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_4_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29713),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29694),
            .ce(),
            .sr(N__46969));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_12_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_12_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_12_5_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_12_5_3  (
            .in0(N__29682),
            .in1(N__29636),
            .in2(_gnd_net_),
            .in3(N__41168),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47509),
            .ce(N__32029),
            .sr(N__46976));
    defparam \phase_controller_inst1.start_timer_hc_LC_12_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_6_0 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_12_6_0  (
            .in0(N__46466),
            .in1(N__30153),
            .in2(N__33131),
            .in3(N__29613),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47496),
            .ce(),
            .sr(N__46982));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_12_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_12_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_12_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_12_6_1  (
            .in0(N__30152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47496),
            .ce(),
            .sr(N__46982));
    defparam \phase_controller_inst1.stoper_hc.running_LC_12_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_12_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_12_6_2 .LUT_INIT=16'b1101111100001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_12_6_2  (
            .in0(N__32158),
            .in1(N__30758),
            .in2(N__30137),
            .in3(N__29589),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47496),
            .ce(),
            .sr(N__46982));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__32157),
            .in2(_gnd_net_),
            .in3(N__32137),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_12_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_12_6_4 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_12_6_4  (
            .in0(N__30128),
            .in1(N__29588),
            .in2(_gnd_net_),
            .in3(N__30150),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_6_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30162),
            .in3(N__32138),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_6 .LUT_INIT=16'b1100010011100100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_6  (
            .in0(N__32159),
            .in1(N__32731),
            .in2(N__30138),
            .in3(N__30759),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47496),
            .ce(),
            .sr(N__46982));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_6_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_6_7  (
            .in0(N__30151),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30129),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_12_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_12_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__30105),
            .in2(N__30093),
            .in3(N__31822),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_12_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_12_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__30084),
            .in2(N__30057),
            .in3(N__30072),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_12_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_12_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__30048),
            .in2(N__30015),
            .in3(N__30036),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_12_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_12_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__30006),
            .in2(N__29979),
            .in3(N__29994),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_12_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_12_7_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_12_7_4  (
            .in0(N__29970),
            .in1(N__29955),
            .in2(N__29946),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_12_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_12_7_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_12_7_5  (
            .in0(N__30429),
            .in1(N__30414),
            .in2(N__30402),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_12_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_12_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(N__30390),
            .in2(N__30366),
            .in3(N__30381),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_12_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_12_7_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_12_7_7  (
            .in0(N__30357),
            .in1(N__30342),
            .in2(N__30324),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_12_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_12_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__30312),
            .in2(N__30282),
            .in3(N__30300),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_12_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_12_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__30273),
            .in2(N__30246),
            .in3(N__30261),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_12_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_12_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__30237),
            .in2(N__30207),
            .in3(N__30225),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_12_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_12_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__30195),
            .in2(N__30171),
            .in3(N__30186),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_12_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_12_8_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_12_8_4  (
            .in0(N__30666),
            .in1(N__30651),
            .in2(N__30636),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_12_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_12_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_12_8_5  (
            .in0(N__30624),
            .in1(N__30594),
            .in2(N__30606),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_12_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_12_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__30588),
            .in2(N__30564),
            .in3(N__30579),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_12_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_12_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__30555),
            .in2(N__30546),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_12_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__30531),
            .in2(N__30519),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_12_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_12_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__30504),
            .in2(N__30495),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_12_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_12_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__30483),
            .in2(N__30471),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_12_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_12_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__30456),
            .in2(N__30444),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_12_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_12_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__30846),
            .in2(N__30834),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_12_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_12_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__30819),
            .in2(N__30807),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__30792),
            .in2(N__30786),
            .in3(N__30765),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30762),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__30747),
            .in2(N__30741),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_10_1  (
            .in0(N__32455),
            .in1(N__30720),
            .in2(_gnd_net_),
            .in3(N__30708),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__47453),
            .ce(),
            .sr(N__47012));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_10_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_10_2  (
            .in0(N__32459),
            .in1(N__30696),
            .in2(N__30705),
            .in3(N__30684),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__47453),
            .ce(),
            .sr(N__47012));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_10_3  (
            .in0(N__32456),
            .in1(N__30681),
            .in2(_gnd_net_),
            .in3(N__30669),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__47453),
            .ce(),
            .sr(N__47012));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_10_4  (
            .in0(N__32460),
            .in1(N__30966),
            .in2(_gnd_net_),
            .in3(N__30954),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__47453),
            .ce(),
            .sr(N__47012));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_10_5  (
            .in0(N__32457),
            .in1(N__30951),
            .in2(_gnd_net_),
            .in3(N__30939),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__47453),
            .ce(),
            .sr(N__47012));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_10_6  (
            .in0(N__32461),
            .in1(N__30936),
            .in2(_gnd_net_),
            .in3(N__30924),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__47453),
            .ce(),
            .sr(N__47012));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_10_7  (
            .in0(N__32458),
            .in1(N__30921),
            .in2(_gnd_net_),
            .in3(N__30909),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__47453),
            .ce(),
            .sr(N__47012));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_11_0  (
            .in0(N__32450),
            .in1(N__30906),
            .in2(_gnd_net_),
            .in3(N__30894),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__47443),
            .ce(),
            .sr(N__47019));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_11_1  (
            .in0(N__32462),
            .in1(N__30891),
            .in2(_gnd_net_),
            .in3(N__30879),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__47443),
            .ce(),
            .sr(N__47019));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_11_2  (
            .in0(N__32447),
            .in1(N__30876),
            .in2(_gnd_net_),
            .in3(N__30864),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__47443),
            .ce(),
            .sr(N__47019));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_11_3  (
            .in0(N__32463),
            .in1(N__30861),
            .in2(_gnd_net_),
            .in3(N__30849),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__47443),
            .ce(),
            .sr(N__47019));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_11_4  (
            .in0(N__32448),
            .in1(N__31161),
            .in2(_gnd_net_),
            .in3(N__31149),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__47443),
            .ce(),
            .sr(N__47019));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_11_5  (
            .in0(N__32464),
            .in1(N__31146),
            .in2(_gnd_net_),
            .in3(N__31134),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__47443),
            .ce(),
            .sr(N__47019));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_11_6  (
            .in0(N__32449),
            .in1(N__31131),
            .in2(_gnd_net_),
            .in3(N__31119),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__47443),
            .ce(),
            .sr(N__47019));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_11_7  (
            .in0(N__32465),
            .in1(N__31106),
            .in2(_gnd_net_),
            .in3(N__31092),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__47443),
            .ce(),
            .sr(N__47019));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_12_0  (
            .in0(N__32451),
            .in1(N__31087),
            .in2(_gnd_net_),
            .in3(N__31071),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__47438),
            .ce(),
            .sr(N__47026));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_12_1  (
            .in0(N__32466),
            .in1(N__31061),
            .in2(_gnd_net_),
            .in3(N__31047),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__47438),
            .ce(),
            .sr(N__47026));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_12_2  (
            .in0(N__32452),
            .in1(N__31034),
            .in2(_gnd_net_),
            .in3(N__31020),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__47438),
            .ce(),
            .sr(N__47026));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_12_3  (
            .in0(N__32467),
            .in1(N__31010),
            .in2(_gnd_net_),
            .in3(N__30996),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__47438),
            .ce(),
            .sr(N__47026));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_12_4  (
            .in0(N__32453),
            .in1(N__30983),
            .in2(_gnd_net_),
            .in3(N__30969),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__47438),
            .ce(),
            .sr(N__47026));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_12_5  (
            .in0(N__32468),
            .in1(N__31364),
            .in2(_gnd_net_),
            .in3(N__31350),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__47438),
            .ce(),
            .sr(N__47026));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_12_6  (
            .in0(N__32454),
            .in1(N__31340),
            .in2(_gnd_net_),
            .in3(N__31326),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__47438),
            .ce(),
            .sr(N__47026));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_12_7  (
            .in0(N__32469),
            .in1(N__31313),
            .in2(_gnd_net_),
            .in3(N__31299),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__47438),
            .ce(),
            .sr(N__47026));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_13_0  (
            .in0(N__32474),
            .in1(N__31294),
            .in2(_gnd_net_),
            .in3(N__31278),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__47433),
            .ce(),
            .sr(N__47032));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_13_1  (
            .in0(N__32478),
            .in1(N__31267),
            .in2(_gnd_net_),
            .in3(N__31248),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__47433),
            .ce(),
            .sr(N__47032));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_13_2  (
            .in0(N__32475),
            .in1(N__31237),
            .in2(_gnd_net_),
            .in3(N__31215),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__47433),
            .ce(),
            .sr(N__47032));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_13_3  (
            .in0(N__32479),
            .in1(N__31202),
            .in2(_gnd_net_),
            .in3(N__31188),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__47433),
            .ce(),
            .sr(N__47032));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_13_4  (
            .in0(N__32476),
            .in1(N__31178),
            .in2(_gnd_net_),
            .in3(N__31164),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__47433),
            .ce(),
            .sr(N__47032));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_13_5  (
            .in0(N__32480),
            .in1(N__31491),
            .in2(_gnd_net_),
            .in3(N__31473),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__47433),
            .ce(),
            .sr(N__47032));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_13_6  (
            .in0(N__32477),
            .in1(N__31451),
            .in2(_gnd_net_),
            .in3(N__31470),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47433),
            .ce(),
            .sr(N__47032));
    defparam \phase_controller_inst1.state_2_LC_12_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_12_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_12_14_5 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst1.state_2_LC_12_14_5  (
            .in0(N__32714),
            .in1(N__31759),
            .in2(N__32754),
            .in3(N__31436),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47429),
            .ce(),
            .sr(N__47038));
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_12_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_12_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNIE87F_2_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__32713),
            .in2(_gnd_net_),
            .in3(N__32749),
            .lcout(\phase_controller_inst1.state_RNIE87FZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6  (
            .in0(N__40580),
            .in1(N__42487),
            .in2(N__40230),
            .in3(N__36848),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_16_0 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_16_0  (
            .in0(N__39954),
            .in1(N__40576),
            .in2(N__37034),
            .in3(N__42621),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_12_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_12_16_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_12_16_1  (
            .in0(N__40573),
            .in1(N__39956),
            .in2(N__42453),
            .in3(N__36816),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_16_2 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_16_2  (
            .in0(N__37472),
            .in1(N__40571),
            .in2(N__32807),
            .in3(N__39498),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_12_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_12_16_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_12_16_3  (
            .in0(N__40575),
            .in1(N__39958),
            .in2(N__42851),
            .in3(N__37163),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_12_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_12_16_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_12_16_6  (
            .in0(N__39955),
            .in1(N__40572),
            .in2(N__42495),
            .in3(N__36849),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_16_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_16_7  (
            .in0(N__40574),
            .in1(N__39957),
            .in2(N__42360),
            .in3(N__37196),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__32921),
            .in2(N__32892),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__32796),
            .in2(N__32775),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__32625),
            .in2(N__39965),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__39791),
            .in2(N__31503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__32847),
            .in2(N__39966),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__39795),
            .in2(N__32841),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(N__32832),
            .in2(N__39967),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__39799),
            .in2(N__31524),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__39803),
            .in2(N__32826),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__32910),
            .in2(N__39968),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__39807),
            .in2(N__32817),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__32982),
            .in2(N__39969),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__39811),
            .in2(N__32871),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__32904),
            .in2(N__39970),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__39815),
            .in2(N__34617),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__32862),
            .in2(N__39971),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__32898),
            .in2(N__40137),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__39995),
            .in2(N__32856),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__32877),
            .in2(N__40138),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__39999),
            .in2(N__34791),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__34671),
            .in2(N__40139),
            .in3(N__31581),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__40003),
            .in2(N__32952),
            .in3(N__31566),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__38088),
            .in2(N__40140),
            .in3(N__31551),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(N__40007),
            .in2(N__37272),
            .in3(N__31536),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__40021),
            .in2(N__37323),
            .in3(N__31527),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__37809),
            .in2(N__40144),
            .in3(N__31668),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__40025),
            .in2(N__39663),
            .in3(N__31656),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__32934),
            .in2(N__40145),
            .in3(N__31641),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__40029),
            .in2(N__32976),
            .in3(N__31629),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__38289),
            .in2(N__40146),
            .in3(N__31617),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__40033),
            .in2(N__37338),
            .in3(N__31605),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_20_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_20_7  (
            .in0(N__40034),
            .in1(N__40444),
            .in2(_gnd_net_),
            .in3(N__31602),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_LC_12_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_12_21_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_12_21_1  (
            .in0(N__31784),
            .in1(N__31769),
            .in2(N__33024),
            .in3(N__33041),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47419),
            .ce(),
            .sr(N__47065));
    defparam \current_shift_inst.timer_s1.running_LC_12_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_12_21_4 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_12_21_4  (
            .in0(N__33042),
            .in1(N__33020),
            .in2(_gnd_net_),
            .in3(N__41306),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47419),
            .ce(),
            .sr(N__47065));
    defparam \phase_controller_inst1.S1_LC_12_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_12_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31770),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47419),
            .ce(),
            .sr(N__47065));
    defparam \current_shift_inst.start_timer_s1_LC_12_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_12_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_12_21_7 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_12_21_7  (
            .in0(N__31783),
            .in1(N__33040),
            .in2(_gnd_net_),
            .in3(N__31768),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47419),
            .ce(),
            .sr(N__47065));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0  (
            .in0(N__35839),
            .in1(N__36078),
            .in2(N__36000),
            .in3(N__31734),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1  (
            .in0(N__36079),
            .in1(N__35840),
            .in2(N__31728),
            .in3(N__35950),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2  (
            .in0(N__35841),
            .in1(N__36080),
            .in2(N__36001),
            .in3(N__31719),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3  (
            .in0(N__36081),
            .in1(N__35951),
            .in2(N__31713),
            .in3(N__35842),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5  (
            .in0(N__36075),
            .in1(N__35939),
            .in2(N__31704),
            .in3(N__35836),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_24_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_24_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_24_6  (
            .in0(N__35838),
            .in1(N__36077),
            .in2(N__35999),
            .in3(N__31695),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7  (
            .in0(N__36076),
            .in1(N__35943),
            .in2(N__31689),
            .in3(N__35837),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_2 .LUT_INIT=16'b1101110111001111;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_2  (
            .in0(N__35852),
            .in1(N__32187),
            .in2(N__36090),
            .in3(N__35953),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_7 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_7  (
            .in0(N__35952),
            .in1(N__35853),
            .in2(N__32181),
            .in3(N__36088),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_4 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_4 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_4  (
            .in0(N__47121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_1_LC_13_3_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_13_3_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_13_3_4 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst2.state_1_LC_13_3_4  (
            .in0(N__35731),
            .in1(N__41927),
            .in2(_gnd_net_),
            .in3(N__35709),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47543),
            .ce(),
            .sr(N__46959));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_4_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_4_2  (
            .in0(N__38180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39576),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_13_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_13_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_13_5_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_31_LC_13_5_3  (
            .in0(N__44706),
            .in1(N__44321),
            .in2(_gnd_net_),
            .in3(N__48332),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47523),
            .ce(N__47825),
            .sr(N__46970));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_6_1 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_6_1  (
            .in0(N__46563),
            .in1(N__36945),
            .in2(N__38854),
            .in3(N__47874),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47512),
            .ce(),
            .sr(N__46977));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_6_2 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_6_2  (
            .in0(N__32160),
            .in1(N__31826),
            .in2(N__32142),
            .in3(N__31984),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47512),
            .ce(),
            .sr(N__46977));
    defparam \phase_controller_inst2.start_timer_hc_LC_13_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_13_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_13_6_3 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_13_6_3  (
            .in0(N__31806),
            .in1(N__46456),
            .in2(N__32295),
            .in3(N__35708),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47512),
            .ce(),
            .sr(N__46977));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_6_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_6_4  (
            .in0(N__32215),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32290),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_13_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_13_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_13_6_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_13_6_5  (
            .in0(N__32294),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47512),
            .ce(),
            .sr(N__46977));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_6_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_6_6  (
            .in0(N__32214),
            .in1(N__32319),
            .in2(_gnd_net_),
            .in3(N__32289),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst2.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_13_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_13_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_13_6_7 .LUT_INIT=16'b1011101000001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_13_6_7  (
            .in0(N__38122),
            .in1(N__32256),
            .in2(N__32232),
            .in3(N__32216),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47512),
            .ce(),
            .sr(N__46977));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_7_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__33380),
            .in2(N__36231),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47498),
            .ce(N__36196),
            .sr(N__46983));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__33353),
            .in2(N__33414),
            .in3(N__32199),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47498),
            .ce(N__36196),
            .sr(N__46983));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__33332),
            .in2(N__33384),
            .in3(N__32196),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47498),
            .ce(N__36196),
            .sr(N__46983));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__33354),
            .in2(N__33719),
            .in3(N__32193),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47498),
            .ce(N__36196),
            .sr(N__46983));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__33333),
            .in2(N__33692),
            .in3(N__32190),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47498),
            .ce(N__36196),
            .sr(N__46983));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__33659),
            .in2(N__33720),
            .in3(N__32514),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47498),
            .ce(N__36196),
            .sr(N__46983));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(N__33625),
            .in2(N__33693),
            .in3(N__32511),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47498),
            .ce(N__36196),
            .sr(N__46983));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__33595),
            .in2(N__33663),
            .in3(N__32508),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47498),
            .ce(N__36196),
            .sr(N__46983));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(N__33633),
            .in2(N__33575),
            .in3(N__32505),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47486),
            .ce(N__36195),
            .sr(N__46990));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__33548),
            .in2(N__33606),
            .in3(N__32502),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47486),
            .ce(N__36195),
            .sr(N__46990));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__33527),
            .in2(N__33576),
            .in3(N__32499),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47486),
            .ce(N__36195),
            .sr(N__46990));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__33549),
            .in2(N__33938),
            .in3(N__32496),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47486),
            .ce(N__36195),
            .sr(N__46990));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(N__33528),
            .in2(N__33911),
            .in3(N__32493),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47486),
            .ce(N__36195),
            .sr(N__46990));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__33881),
            .in2(N__33939),
            .in3(N__32490),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47486),
            .ce(N__36195),
            .sr(N__46990));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__33844),
            .in2(N__33912),
            .in3(N__32541),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47486),
            .ce(N__36195),
            .sr(N__46990));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__33814),
            .in2(N__33882),
            .in3(N__32538),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47486),
            .ce(N__36195),
            .sr(N__46990));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__33794),
            .in2(N__33852),
            .in3(N__32535),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47473),
            .ce(N__36194),
            .sr(N__46999));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__33770),
            .in2(N__33825),
            .in3(N__32532),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47473),
            .ce(N__36194),
            .sr(N__46999));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__33795),
            .in2(N__33749),
            .in3(N__32529),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47473),
            .ce(N__36194),
            .sr(N__46999));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__33771),
            .in2(N__34217),
            .in3(N__32526),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47473),
            .ce(N__36194),
            .sr(N__46999));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__34190),
            .in2(N__33750),
            .in3(N__32523),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47473),
            .ce(N__36194),
            .sr(N__46999));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__34169),
            .in2(N__34218),
            .in3(N__32520),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47473),
            .ce(N__36194),
            .sr(N__46999));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__34191),
            .in2(N__34139),
            .in3(N__32517),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47473),
            .ce(N__36194),
            .sr(N__46999));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__34099),
            .in2(N__34170),
            .in3(N__32562),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47473),
            .ce(N__36194),
            .sr(N__46999));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__34140),
            .in2(N__34079),
            .in3(N__32559),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47463),
            .ce(N__36178),
            .sr(N__47007));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__34052),
            .in2(N__34110),
            .in3(N__32556),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47463),
            .ce(N__36178),
            .sr(N__47007));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__34032),
            .in2(N__34080),
            .in3(N__32553),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47463),
            .ce(N__36178),
            .sr(N__47007));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__34053),
            .in2(N__34011),
            .in3(N__32550),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47463),
            .ce(N__36178),
            .sr(N__47007));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32547),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47463),
            .ce(N__36178),
            .sr(N__47007));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_13_11_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_13_11_0  (
            .in0(N__39066),
            .in1(N__39089),
            .in2(N__32619),
            .in3(N__32604),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_11_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_11_1  (
            .in0(N__32603),
            .in1(N__39065),
            .in2(N__39093),
            .in3(N__32615),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_13_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_13_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_13_11_2  (
            .in0(N__36292),
            .in1(N__36305),
            .in2(_gnd_net_),
            .in3(N__48263),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(elapsed_time_ns_1_RNI1CPBB_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_13_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_13_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_13_11_3 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_23_LC_13_11_3  (
            .in0(N__48266),
            .in1(N__36293),
            .in2(N__32544),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47455),
            .ce(N__47875),
            .sr(N__47013));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_13_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_13_11_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_13_11_4  (
            .in0(N__36369),
            .in1(N__48264),
            .in2(_gnd_net_),
            .in3(N__36332),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_13_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_13_11_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_22_LC_13_11_5  (
            .in0(N__48265),
            .in1(_gnd_net_),
            .in2(N__32607),
            .in3(N__36370),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47455),
            .ce(N__47875),
            .sr(N__47013));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_13_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_13_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_13_11_6  (
            .in0(N__45340),
            .in1(N__45378),
            .in2(_gnd_net_),
            .in3(N__48267),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47455),
            .ce(N__47875),
            .sr(N__47013));
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_13_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_13_12_0 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_13_12_0  (
            .in0(N__32590),
            .in1(N__39232),
            .in2(N__39272),
            .in3(N__32578),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_13_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_13_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_13_12_1  (
            .in0(N__48333),
            .in1(N__41833),
            .in2(_gnd_net_),
            .in3(N__41798),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_13_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_13_12_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_30_LC_13_12_2  (
            .in0(N__41834),
            .in1(_gnd_net_),
            .in2(N__32595),
            .in3(N__48335),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47445),
            .ce(N__47877),
            .sr(N__47020));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_12_3 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_12_3  (
            .in0(N__32580),
            .in1(N__32592),
            .in2(N__39237),
            .in3(N__39271),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_13_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_13_12_6 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_13_12_6  (
            .in0(N__32591),
            .in1(N__39233),
            .in2(N__39273),
            .in3(N__32579),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_13_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_13_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_13_12_7  (
            .in0(N__48334),
            .in1(N__46172),
            .in2(_gnd_net_),
            .in3(N__46146),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47445),
            .ce(N__47877),
            .sr(N__47020));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33078),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43170),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__43229),
            .sr(N__47027));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_6  (
            .in0(N__43200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__43229),
            .sr(N__47027));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_1  (
            .in0(N__38005),
            .in1(N__36912),
            .in2(_gnd_net_),
            .in3(N__33079),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42576),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_14_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_14_7  (
            .in0(N__33155),
            .in1(N__33461),
            .in2(N__32753),
            .in3(N__32715),
            .lcout(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_13_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_13_15_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_13_15_1  (
            .in0(N__32654),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46433),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_5 .LUT_INIT=16'b1101000011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_5  (
            .in0(N__47576),
            .in1(N__32689),
            .in2(N__46656),
            .in3(N__46546),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47431),
            .ce(),
            .sr(N__47039));
    defparam \phase_controller_inst1.state_4_LC_13_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_13_15_6 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_13_15_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.state_4_LC_13_15_6  (
            .in0(N__46434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32653),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47431),
            .ce(),
            .sr(N__47039));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_16_2  (
            .in0(N__40577),
            .in1(N__46271),
            .in2(N__40231),
            .in3(N__36881),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_13_16_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_13_16_3  (
            .in0(N__36815),
            .in1(N__40578),
            .in2(N__40232),
            .in3(N__42449),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_16_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_16_4  (
            .in0(N__38006),
            .in1(N__42488),
            .in2(_gnd_net_),
            .in3(N__36847),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_16_7 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_16_7  (
            .in0(N__42399),
            .in1(N__40150),
            .in2(N__37548),
            .in3(N__40579),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_13_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_13_17_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_13_17_0  (
            .in0(N__40483),
            .in1(N__40112),
            .in2(N__42359),
            .in3(N__37197),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_13_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_13_17_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_13_17_1  (
            .in0(N__40113),
            .in1(N__40484),
            .in2(N__37584),
            .in3(N__42800),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_17_2 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_17_2  (
            .in0(N__40486),
            .in1(N__37104),
            .in2(N__42714),
            .in3(N__40111),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_17_3  (
            .in0(N__38016),
            .in1(N__42445),
            .in2(_gnd_net_),
            .in3(N__36814),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_4  (
            .in0(N__40482),
            .in1(N__37473),
            .in2(N__32808),
            .in3(N__39497),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_17_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_17_5  (
            .in0(N__35507),
            .in1(N__32766),
            .in2(_gnd_net_),
            .in3(N__34757),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_17_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_17_6  (
            .in0(N__32891),
            .in1(_gnd_net_),
            .in2(N__32928),
            .in3(N__35508),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_17_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_17_7  (
            .in0(N__40114),
            .in1(N__40485),
            .in2(N__42756),
            .in3(N__37130),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_18_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_18_0  (
            .in0(N__40448),
            .in1(N__40200),
            .in2(N__37038),
            .in3(N__42620),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_18_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_18_1  (
            .in0(N__40202),
            .in1(N__40450),
            .in2(N__37782),
            .in3(N__43088),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_18_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_18_2  (
            .in0(N__40445),
            .in1(N__33096),
            .in2(_gnd_net_),
            .in3(N__33087),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_3  (
            .in0(N__40204),
            .in1(N__40452),
            .in2(N__37623),
            .in3(N__43007),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_18_4 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_18_4  (
            .in0(N__40447),
            .in1(N__40199),
            .in2(N__37074),
            .in3(N__42671),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_18_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_18_5  (
            .in0(N__40201),
            .in1(N__40449),
            .in2(N__43140),
            .in3(N__37380),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_13_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_13_18_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_13_18_6  (
            .in0(N__40451),
            .in1(N__40203),
            .in2(N__43050),
            .in3(N__37716),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_18_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_18_7  (
            .in0(N__40198),
            .in1(N__40446),
            .in2(N__46377),
            .in3(N__37434),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_19_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_19_1  (
            .in0(N__40196),
            .in1(N__40442),
            .in2(N__37881),
            .in3(N__43320),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_19_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_19_3  (
            .in0(N__40195),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40443),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5  (
            .in0(N__40197),
            .in1(N__40441),
            .in2(N__37239),
            .in3(N__42893),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6  (
            .in0(N__37957),
            .in1(N__42892),
            .in2(_gnd_net_),
            .in3(N__37235),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7  (
            .in0(N__43192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47425),
            .ce(N__43227),
            .sr(N__47058));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_20_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_20_1  (
            .in0(N__40362),
            .in1(N__43352),
            .in2(N__40256),
            .in3(N__38072),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_20_2 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_20_2  (
            .in0(N__43353),
            .in1(N__40363),
            .in2(N__38073),
            .in3(N__40208),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43193),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47422),
            .ce(N__43226),
            .sr(N__47061));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36924),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_20_6 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_20_6  (
            .in0(N__33086),
            .in1(N__40361),
            .in2(N__33060),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_2 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_2  (
            .in0(N__41302),
            .in1(N__33019),
            .in2(_gnd_net_),
            .in3(N__33039),
            .lcout(\current_shift_inst.timer_s1.N_163_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(N__41301),
            .in2(_gnd_net_),
            .in3(N__33018),
            .lcout(\current_shift_inst.timer_s1.N_162_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__35208),
            .in2(_gnd_net_),
            .in3(N__38276),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_200_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_21_6 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_21_6  (
            .in0(N__35209),
            .in1(_gnd_net_),
            .in2(N__38280),
            .in3(N__38255),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_201_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_13_22_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_13_22_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_13_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_13_22_0  (
            .in0(N__34962),
            .in1(N__35102),
            .in2(_gnd_net_),
            .in3(N__32991),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__47421),
            .ce(),
            .sr(N__47066));
    defparam \pwm_generator_inst.counter_1_LC_13_22_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_13_22_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_13_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_13_22_1  (
            .in0(N__34956),
            .in1(N__35036),
            .in2(_gnd_net_),
            .in3(N__32988),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__47421),
            .ce(),
            .sr(N__47066));
    defparam \pwm_generator_inst.counter_2_LC_13_22_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_13_22_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_13_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_13_22_2  (
            .in0(N__34963),
            .in1(N__35123),
            .in2(_gnd_net_),
            .in3(N__32985),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__47421),
            .ce(),
            .sr(N__47066));
    defparam \pwm_generator_inst.counter_3_LC_13_22_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_13_22_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_13_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_13_22_3  (
            .in0(N__34957),
            .in1(N__35060),
            .in2(_gnd_net_),
            .in3(N__33180),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__47421),
            .ce(),
            .sr(N__47066));
    defparam \pwm_generator_inst.counter_4_LC_13_22_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_13_22_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_13_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_13_22_4  (
            .in0(N__34964),
            .in1(N__35081),
            .in2(_gnd_net_),
            .in3(N__33177),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__47421),
            .ce(),
            .sr(N__47066));
    defparam \pwm_generator_inst.counter_5_LC_13_22_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_13_22_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_13_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_13_22_5  (
            .in0(N__34958),
            .in1(N__34984),
            .in2(_gnd_net_),
            .in3(N__33174),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__47421),
            .ce(),
            .sr(N__47066));
    defparam \pwm_generator_inst.counter_6_LC_13_22_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_13_22_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_13_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_13_22_6  (
            .in0(N__34965),
            .in1(N__35008),
            .in2(_gnd_net_),
            .in3(N__33171),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__47421),
            .ce(),
            .sr(N__47066));
    defparam \pwm_generator_inst.counter_7_LC_13_22_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_13_22_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_13_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_13_22_7  (
            .in0(N__34959),
            .in1(N__35144),
            .in2(_gnd_net_),
            .in3(N__33168),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__47421),
            .ce(),
            .sr(N__47066));
    defparam \pwm_generator_inst.counter_8_LC_13_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_13_23_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_13_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_13_23_0  (
            .in0(N__34961),
            .in1(N__35165),
            .in2(_gnd_net_),
            .in3(N__33165),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__47418),
            .ce(),
            .sr(N__47070));
    defparam \pwm_generator_inst.counter_9_LC_13_23_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_13_23_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_13_23_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_13_23_1  (
            .in0(N__35186),
            .in1(N__34960),
            .in2(_gnd_net_),
            .in3(N__33162),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47418),
            .ce(),
            .sr(N__47070));
    defparam \phase_controller_inst1.state_1_LC_13_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_13_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_13_23_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst1.state_1_LC_13_23_3  (
            .in0(N__33159),
            .in1(N__33453),
            .in2(_gnd_net_),
            .in3(N__33132),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47418),
            .ce(),
            .sr(N__47070));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__33102),
            .in2(N__35802),
            .in3(N__35103),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1  (
            .in0(N__35037),
            .in1(N__33303),
            .in2(N__33312),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__33285),
            .in2(N__33297),
            .in3(N__35124),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__33267),
            .in2(N__33279),
            .in3(N__35061),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4  (
            .in0(N__35082),
            .in1(N__33249),
            .in2(N__33261),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__33234),
            .in2(N__33243),
            .in3(N__34986),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6  (
            .in0(N__35010),
            .in1(N__33219),
            .in2(N__33228),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__33204),
            .in2(N__33213),
            .in3(N__35145),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__33186),
            .in2(N__33198),
            .in3(N__35166),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__33498),
            .in2(N__33507),
            .in3(N__35187),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_13_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_13_25_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_13_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33492),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47416),
            .ce(),
            .sr(N__47078));
    defparam \phase_controller_inst1.S2_LC_13_29_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_29_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_29_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_29_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33457),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47412),
            .ce(),
            .sr(N__47092));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_4_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_4_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33407),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47544),
            .ce(N__36204),
            .sr(N__46960));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_5_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_5_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_5_0  (
            .in0(N__34343),
            .in1(N__36220),
            .in2(_gnd_net_),
            .in3(N__33417),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__47533),
            .ce(N__33993),
            .sr(N__46964));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_5_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_5_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_5_1  (
            .in0(N__34347),
            .in1(N__33406),
            .in2(_gnd_net_),
            .in3(N__33387),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__47533),
            .ce(N__33993),
            .sr(N__46964));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_5_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_5_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_5_2  (
            .in0(N__34344),
            .in1(N__33379),
            .in2(_gnd_net_),
            .in3(N__33357),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__47533),
            .ce(N__33993),
            .sr(N__46964));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_5_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_5_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_5_3  (
            .in0(N__34348),
            .in1(N__33352),
            .in2(_gnd_net_),
            .in3(N__33336),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__47533),
            .ce(N__33993),
            .sr(N__46964));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_5_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_5_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_5_4  (
            .in0(N__34345),
            .in1(N__33331),
            .in2(_gnd_net_),
            .in3(N__33315),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__47533),
            .ce(N__33993),
            .sr(N__46964));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_5_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_5_5  (
            .in0(N__34349),
            .in1(N__33712),
            .in2(_gnd_net_),
            .in3(N__33696),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__47533),
            .ce(N__33993),
            .sr(N__46964));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_5_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_5_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_5_6  (
            .in0(N__34346),
            .in1(N__33680),
            .in2(_gnd_net_),
            .in3(N__33666),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__47533),
            .ce(N__33993),
            .sr(N__46964));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_5_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_5_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_5_7  (
            .in0(N__34350),
            .in1(N__33652),
            .in2(_gnd_net_),
            .in3(N__33636),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__47533),
            .ce(N__33993),
            .sr(N__46964));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_6_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_6_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_6_0  (
            .in0(N__34342),
            .in1(N__33626),
            .in2(_gnd_net_),
            .in3(N__33609),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__47524),
            .ce(N__33992),
            .sr(N__46971));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_6_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_6_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_6_1  (
            .in0(N__34338),
            .in1(N__33599),
            .in2(_gnd_net_),
            .in3(N__33579),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__47524),
            .ce(N__33992),
            .sr(N__46971));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_6_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_6_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_6_2  (
            .in0(N__34339),
            .in1(N__33568),
            .in2(_gnd_net_),
            .in3(N__33552),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__47524),
            .ce(N__33992),
            .sr(N__46971));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_6_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_6_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_6_3  (
            .in0(N__34335),
            .in1(N__33547),
            .in2(_gnd_net_),
            .in3(N__33531),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__47524),
            .ce(N__33992),
            .sr(N__46971));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_6_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_6_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_6_4  (
            .in0(N__34340),
            .in1(N__33526),
            .in2(_gnd_net_),
            .in3(N__33510),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__47524),
            .ce(N__33992),
            .sr(N__46971));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_6_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_6_5  (
            .in0(N__34336),
            .in1(N__33931),
            .in2(_gnd_net_),
            .in3(N__33915),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__47524),
            .ce(N__33992),
            .sr(N__46971));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_6_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_6_6  (
            .in0(N__34341),
            .in1(N__33899),
            .in2(_gnd_net_),
            .in3(N__33885),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__47524),
            .ce(N__33992),
            .sr(N__46971));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_6_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_6_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_6_7  (
            .in0(N__34337),
            .in1(N__33874),
            .in2(_gnd_net_),
            .in3(N__33855),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__47524),
            .ce(N__33992),
            .sr(N__46971));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_7_0  (
            .in0(N__34307),
            .in1(N__33845),
            .in2(_gnd_net_),
            .in3(N__33828),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__47513),
            .ce(N__33991),
            .sr(N__46978));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_7_1  (
            .in0(N__34331),
            .in1(N__33818),
            .in2(_gnd_net_),
            .in3(N__33798),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__47513),
            .ce(N__33991),
            .sr(N__46978));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_7_2  (
            .in0(N__34308),
            .in1(N__33793),
            .in2(_gnd_net_),
            .in3(N__33774),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__47513),
            .ce(N__33991),
            .sr(N__46978));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_7_3  (
            .in0(N__34332),
            .in1(N__33769),
            .in2(_gnd_net_),
            .in3(N__33753),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__47513),
            .ce(N__33991),
            .sr(N__46978));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_7_4  (
            .in0(N__34309),
            .in1(N__33737),
            .in2(_gnd_net_),
            .in3(N__33723),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__47513),
            .ce(N__33991),
            .sr(N__46978));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_7_5  (
            .in0(N__34333),
            .in1(N__34210),
            .in2(_gnd_net_),
            .in3(N__34194),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__47513),
            .ce(N__33991),
            .sr(N__46978));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_7_6  (
            .in0(N__34310),
            .in1(N__34189),
            .in2(_gnd_net_),
            .in3(N__34173),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__47513),
            .ce(N__33991),
            .sr(N__46978));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_7_7  (
            .in0(N__34334),
            .in1(N__34162),
            .in2(_gnd_net_),
            .in3(N__34143),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__47513),
            .ce(N__33991),
            .sr(N__46978));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_8_0  (
            .in0(N__34303),
            .in1(N__34135),
            .in2(_gnd_net_),
            .in3(N__34113),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__47499),
            .ce(N__33984),
            .sr(N__46984));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_8_1  (
            .in0(N__34311),
            .in1(N__34103),
            .in2(_gnd_net_),
            .in3(N__34083),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__47499),
            .ce(N__33984),
            .sr(N__46984));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_8_2  (
            .in0(N__34304),
            .in1(N__34072),
            .in2(_gnd_net_),
            .in3(N__34056),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__47499),
            .ce(N__33984),
            .sr(N__46984));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_8_3  (
            .in0(N__34312),
            .in1(N__34051),
            .in2(_gnd_net_),
            .in3(N__34035),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__47499),
            .ce(N__33984),
            .sr(N__46984));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_8_4  (
            .in0(N__34305),
            .in1(N__34031),
            .in2(_gnd_net_),
            .in3(N__34017),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__47499),
            .ce(N__33984),
            .sr(N__46984));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_8_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_8_5  (
            .in0(N__34007),
            .in1(N__34306),
            .in2(_gnd_net_),
            .in3(N__34014),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47499),
            .ce(N__33984),
            .sr(N__46984));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35214),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_14_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_14_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_14_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_14_9_0  (
            .in0(N__48288),
            .in1(N__48426),
            .in2(_gnd_net_),
            .in3(N__48463),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47487),
            .ce(N__47861),
            .sr(N__46991));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_14_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_14_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_14_9_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_14_9_3  (
            .in0(N__45015),
            .in1(N__48291),
            .in2(_gnd_net_),
            .in3(N__44983),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47487),
            .ce(N__47861),
            .sr(N__46991));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_14_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_14_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_14_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_14_9_5  (
            .in0(N__44871),
            .in1(N__48292),
            .in2(_gnd_net_),
            .in3(N__36611),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47487),
            .ce(N__47861),
            .sr(N__46991));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_14_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_14_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_14_9_6  (
            .in0(N__48289),
            .in1(N__45084),
            .in2(_gnd_net_),
            .in3(N__45056),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47487),
            .ce(N__47861),
            .sr(N__46991));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_14_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_14_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_14_9_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_14_9_7  (
            .in0(N__44830),
            .in1(N__48290),
            .in2(_gnd_net_),
            .in3(N__36255),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47487),
            .ce(N__47861),
            .sr(N__46991));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_14_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_14_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_14_10_0  (
            .in0(N__42277),
            .in1(N__41698),
            .in2(N__46147),
            .in3(N__36652),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_14_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_14_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_14_10_1  (
            .in0(N__34224),
            .in1(N__34401),
            .in2(N__34227),
            .in3(N__34407),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_14_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_14_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_14_10_2  (
            .in0(N__48358),
            .in1(N__45520),
            .in2(N__45767),
            .in3(N__41832),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_14_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_14_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_14_10_3  (
            .in0(N__36736),
            .in1(N__45301),
            .in2(N__44286),
            .in3(N__45181),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_10_4  (
            .in0(N__46487),
            .in1(N__36283),
            .in2(N__36375),
            .in3(N__45132),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_14_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_14_10_5 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_14_10_5  (
            .in0(N__45133),
            .in1(N__48336),
            .in2(N__45116),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(elapsed_time_ns_1_RNIV9PBB_0_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_14_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_14_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_14_10_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_21_LC_14_10_6  (
            .in0(N__48337),
            .in1(_gnd_net_),
            .in2(N__34395),
            .in3(N__45134),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47474),
            .ce(N__47876),
            .sr(N__47000));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_14_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_14_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__36495),
            .in2(N__34392),
            .in3(N__38855),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_14_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_14_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__34383),
            .in2(N__36438),
            .in3(N__38823),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_14_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_14_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(N__36381),
            .in2(N__34377),
            .in3(N__38793),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_14_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_14_11_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_14_11_3  (
            .in0(N__38772),
            .in1(N__44586),
            .in2(N__34368),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_14_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_14_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__35688),
            .in2(N__34359),
            .in3(N__38754),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_14_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_14_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__36243),
            .in2(N__34548),
            .in3(N__38736),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_14_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_14_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_14_11_6  (
            .in0(N__39042),
            .in1(N__34536),
            .in2(N__34527),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_14_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_14_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__34518),
            .in2(N__34506),
            .in3(N__39024),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_14_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_14_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__34497),
            .in2(N__34488),
            .in3(N__39006),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_14_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_14_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__34467),
            .in2(N__34479),
            .in3(N__38988),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_14_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_14_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__34461),
            .in2(N__34452),
            .in3(N__38970),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_14_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_14_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__34440),
            .in2(N__34431),
            .in3(N__38952),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_14_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_14_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_14_12_4  (
            .in0(N__38934),
            .in1(N__34413),
            .in2(N__34422),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_14_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_14_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_14_12_5  (
            .in0(N__38916),
            .in1(N__36762),
            .in2(N__34587),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_14_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_14_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__42252),
            .in2(N__34578),
            .in3(N__39210),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_14_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_14_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(N__36708),
            .in2(N__36690),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_14_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_14_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__42174),
            .in2(N__42318),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_14_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_14_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__36549),
            .in2(N__36588),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_14_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_14_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__34569),
            .in2(N__34560),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_14_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_14_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__45819),
            .in2(N__45882),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_14_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_14_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__42162),
            .in2(N__45894),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_14_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_14_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__46053),
            .in2(N__45990),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__34644),
            .in2(N__36984),
            .in3(N__34638),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34635),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42345),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_14_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_14_14_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_14_14_1  (
            .in0(N__38002),
            .in1(N__46267),
            .in2(_gnd_net_),
            .in3(N__36868),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_14_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_14_14_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_14_14_2  (
            .in0(N__42838),
            .in1(N__38004),
            .in2(_gnd_net_),
            .in3(N__37151),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_14_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_14_3  (
            .in0(N__40598),
            .in1(N__40265),
            .in2(N__42801),
            .in3(N__37573),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_14_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_14_14_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_14_14_4  (
            .in0(N__40264),
            .in1(N__40600),
            .in2(N__37500),
            .in3(N__42577),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_14_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_14_5  (
            .in0(N__40599),
            .in1(N__40263),
            .in2(N__42582),
            .in3(N__37498),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_14_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_14_6  (
            .in0(N__42346),
            .in1(N__38003),
            .in2(_gnd_net_),
            .in3(N__37183),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_15_0 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_15_0  (
            .in0(N__42710),
            .in1(N__40601),
            .in2(N__37100),
            .in3(N__40260),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_15_1  (
            .in0(N__38007),
            .in1(N__42709),
            .in2(_gnd_net_),
            .in3(N__37093),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_15_2 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_15_2  (
            .in0(N__37774),
            .in1(N__40261),
            .in2(N__43095),
            .in3(N__40602),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_15_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_15_3  (
            .in0(N__40604),
            .in1(N__46319),
            .in2(N__40272),
            .in3(N__37681),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_15_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_15_4  (
            .in0(N__42670),
            .in1(N__38009),
            .in2(_gnd_net_),
            .in3(N__37054),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_15_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_15_5  (
            .in0(N__38010),
            .in1(N__42613),
            .in2(_gnd_net_),
            .in3(N__37015),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_15_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_15_6  (
            .in0(N__37615),
            .in1(N__40262),
            .in2(N__43008),
            .in3(N__40603),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_15_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_15_7  (
            .in0(N__38008),
            .in1(N__37118),
            .in2(_gnd_net_),
            .in3(N__42742),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_14_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_14_16_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_14_16_0  (
            .in0(N__42933),
            .in1(N__40615),
            .in2(N__40237),
            .in3(N__37654),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_16_1  (
            .in0(N__40617),
            .in1(N__43472),
            .in2(N__40234),
            .in3(N__37915),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_2  (
            .in0(N__43042),
            .in1(N__40612),
            .in2(N__40238),
            .in3(N__37708),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_14_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_14_16_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_14_16_3  (
            .in0(N__40613),
            .in1(N__42965),
            .in2(N__40235),
            .in3(N__37741),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_16_4 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_16_4  (
            .in0(N__37234),
            .in1(N__42894),
            .in2(N__40236),
            .in3(N__40616),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_14_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_14_16_5 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_14_16_5  (
            .in0(N__43428),
            .in1(N__40170),
            .in2(N__40628),
            .in3(N__37828),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_14_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_14_16_6 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_14_16_6  (
            .in0(N__42966),
            .in1(N__40614),
            .in2(N__37743),
            .in3(N__40163),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_16_7  (
            .in0(N__40621),
            .in1(N__43319),
            .in2(N__40233),
            .in3(N__37873),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_14_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__39437),
            .in2(N__34761),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_14_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__35525),
            .in2(N__37443),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_14_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__34737),
            .in2(N__35588),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_14_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__35529),
            .in2(N__34896),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_14_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_14_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__34887),
            .in2(N__35589),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_14_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_14_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__35533),
            .in2(N__37515),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_14_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_14_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__34881),
            .in2(N__35590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_14_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_14_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__35537),
            .in2(N__34872),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_14_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__37554),
            .in2(N__35587),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_14_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_14_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__35524),
            .in2(N__34860),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_14_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_14_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__34848),
            .in2(N__35584),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_14_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_14_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__35512),
            .in2(N__37404),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_14_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_14_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__34917),
            .in2(N__35585),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_14_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_14_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__35516),
            .in2(N__34908),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_14_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_14_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__37479),
            .in2(N__35586),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_14_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_14_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__35520),
            .in2(N__37347),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_14_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_14_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__35414),
            .in2(N__37752),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_14_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_14_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__37689),
            .in2(N__35503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_14_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_14_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__35418),
            .in2(N__37593),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_14_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_14_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__37722),
            .in2(N__35504),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_14_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_14_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__35422),
            .in2(N__37632),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_14_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_14_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__34926),
            .in2(N__35505),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_14_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_14_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__35426),
            .in2(N__37791),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_14_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_14_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__37662),
            .in2(N__35506),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_14_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_14_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__35401),
            .in2(N__37896),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_14_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_14_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__37887),
            .in2(N__35500),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_14_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_14_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__35405),
            .in2(N__37845),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_14_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_14_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__38046),
            .in2(N__35501),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_14_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_14_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__35409),
            .in2(N__37854),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_14_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_14_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__38079),
            .in2(N__35502),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_14_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_14_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__35413),
            .in2(N__37800),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_14_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_14_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__40570),
            .in2(_gnd_net_),
            .in3(N__35301),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_14_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_14_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_14_21_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_14_21_4  (
            .in0(N__35210),
            .in1(N__38270),
            .in2(_gnd_net_),
            .in3(N__38256),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47423),
            .ce(),
            .sr(N__47062));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_14_22_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_14_22_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_14_22_3  (
            .in0(N__35182),
            .in1(N__35161),
            .in2(_gnd_net_),
            .in3(N__35143),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_14_22_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_14_22_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__35119),
            .in2(_gnd_net_),
            .in3(N__35098),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_14_22_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_14_22_5 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_14_22_5  (
            .in0(N__35080),
            .in1(N__35059),
            .in2(N__35040),
            .in3(N__35035),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_14_22_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_14_22_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_14_22_6  (
            .in0(N__35016),
            .in1(N__35009),
            .in2(N__34989),
            .in3(N__34985),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_24_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_24_6 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_24_6  (
            .in0(N__36099),
            .in1(N__36089),
            .in2(N__35998),
            .in3(N__35846),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_15_4_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_15_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_15_4_1 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst2.state_0_LC_15_4_1  (
            .in0(N__38106),
            .in1(N__35738),
            .in2(N__41951),
            .in3(N__38214),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47549),
            .ce(),
            .sr(N__46956));
    defparam \phase_controller_inst2.state_3_LC_15_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_15_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_15_4_4 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \phase_controller_inst2.state_3_LC_15_4_4  (
            .in0(N__38181),
            .in1(N__35790),
            .in2(N__39583),
            .in3(N__38198),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47549),
            .ce(),
            .sr(N__46956));
    defparam \phase_controller_inst2.T45_LC_15_4_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.T45_LC_15_4_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T45_LC_15_4_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst2.T45_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(N__35750),
            .in2(_gnd_net_),
            .in3(N__38213),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47549),
            .ce(),
            .sr(N__46956));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_5_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_5_2  (
            .in0(_gnd_net_),
            .in1(N__38362),
            .in2(_gnd_net_),
            .in3(N__38386),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_5_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_5_3  (
            .in0(N__35739),
            .in1(N__41940),
            .in2(N__38456),
            .in3(N__38132),
            .lcout(\phase_controller_inst2.start_timer_tr_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNIG7JF_LC_15_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNIG7JF_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNIG7JF_LC_15_5_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_RNIG7JF_LC_15_5_5  (
            .in0(N__38448),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38131),
            .lcout(\phase_controller_inst2.time_passed_RNIG7JF ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_5_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_5_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_5_7  (
            .in0(N__36604),
            .in1(N__44884),
            .in2(_gnd_net_),
            .in3(N__48268),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_15_6_4  (
            .in0(N__44768),
            .in1(N__44201),
            .in2(_gnd_net_),
            .in3(N__48323),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47534),
            .ce(N__47869),
            .sr(N__46965));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_6_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_15_6_6  (
            .in0(N__44235),
            .in1(N__48324),
            .in2(_gnd_net_),
            .in3(N__44807),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47534),
            .ce(N__47869),
            .sr(N__46965));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_7_0  (
            .in0(N__36399),
            .in1(N__36459),
            .in2(N__44621),
            .in3(N__36513),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_7_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__36230),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47525),
            .ce(N__36203),
            .sr(N__46972));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_7_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_7_4  (
            .in0(N__36539),
            .in1(N__48191),
            .in2(_gnd_net_),
            .in3(N__36514),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_7_5  (
            .in0(N__48190),
            .in1(N__36488),
            .in2(_gnd_net_),
            .in3(N__36460),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_7_6  (
            .in0(N__36400),
            .in1(N__36428),
            .in2(_gnd_net_),
            .in3(N__48192),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_8_0 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_8_0  (
            .in0(N__36120),
            .in1(N__41543),
            .in2(N__36111),
            .in3(N__41522),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_8_1 .LUT_INIT=16'b1101111100001101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_8_1  (
            .in0(N__41544),
            .in1(N__36119),
            .in2(N__41523),
            .in3(N__36107),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_15_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_15_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_15_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_15_8_2  (
            .in0(N__36663),
            .in1(N__48310),
            .in2(_gnd_net_),
            .in3(N__36681),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47514),
            .ce(N__46076),
            .sr(N__46979));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_15_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_15_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_15_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_15_8_3  (
            .in0(N__48307),
            .in1(N__36735),
            .in2(_gnd_net_),
            .in3(N__36756),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47514),
            .ce(N__46076),
            .sr(N__46979));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_15_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_15_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_15_8_4  (
            .in0(N__42283),
            .in1(N__48309),
            .in2(_gnd_net_),
            .in3(N__42303),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47514),
            .ce(N__46076),
            .sr(N__46979));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_15_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_15_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_15_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_15_8_5  (
            .in0(N__48308),
            .in1(N__36535),
            .in2(_gnd_net_),
            .in3(N__36515),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47514),
            .ce(N__46076),
            .sr(N__46979));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_15_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_15_8_6  (
            .in0(N__36484),
            .in1(N__36467),
            .in2(_gnd_net_),
            .in3(N__48314),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47514),
            .ce(N__46076),
            .sr(N__46979));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_15_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_15_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_15_8_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_15_8_7  (
            .in0(N__36407),
            .in1(_gnd_net_),
            .in2(N__48339),
            .in3(N__36424),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47514),
            .ce(N__46076),
            .sr(N__46979));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_9_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_9_0  (
            .in0(N__41657),
            .in1(N__41633),
            .in2(N__36267),
            .in3(N__36321),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_9_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_9_1  (
            .in0(N__36320),
            .in1(N__41658),
            .in2(N__41637),
            .in3(N__36263),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_15_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_15_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_15_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_22_LC_15_9_2  (
            .in0(N__36371),
            .in1(N__48286),
            .in2(_gnd_net_),
            .in3(N__36339),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47500),
            .ce(N__46078),
            .sr(N__46985));
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_15_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_15_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_15_9_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_23_LC_15_9_3  (
            .in0(N__36312),
            .in1(N__48322),
            .in2(_gnd_net_),
            .in3(N__36294),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47500),
            .ce(N__46078),
            .sr(N__46985));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_9_4  (
            .in0(N__44842),
            .in1(N__48284),
            .in2(_gnd_net_),
            .in3(N__36254),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(elapsed_time_ns_1_RNIV8OBB_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_9_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_15_9_5  (
            .in0(N__48285),
            .in1(_gnd_net_),
            .in2(N__36618),
            .in3(N__44843),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47500),
            .ce(N__46078),
            .sr(N__46985));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_15_9_6  (
            .in0(N__36615),
            .in1(N__44885),
            .in2(_gnd_net_),
            .in3(N__48287),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47500),
            .ce(N__46078),
            .sr(N__46985));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_10_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_10_0  (
            .in0(N__39113),
            .in1(N__36557),
            .in2(N__39138),
            .in3(N__36570),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_10_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_10_1  (
            .in0(N__45194),
            .in1(N__48247),
            .in2(_gnd_net_),
            .in3(N__45158),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_15_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_15_10_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_20_LC_15_10_2  (
            .in0(N__48249),
            .in1(_gnd_net_),
            .in2(N__36573),
            .in3(N__45195),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47488),
            .ce(N__47851),
            .sr(N__46992));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_15_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_15_10_3 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_15_10_3  (
            .in0(N__36569),
            .in1(N__39137),
            .in2(N__36561),
            .in3(N__39114),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_15_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_15_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_15_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_15_10_4  (
            .in0(N__48248),
            .in1(N__36540),
            .in2(_gnd_net_),
            .in3(N__36519),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47488),
            .ce(N__47851),
            .sr(N__46992));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_15_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_15_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_15_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_15_10_5  (
            .in0(N__36489),
            .in1(N__36468),
            .in2(_gnd_net_),
            .in3(N__48251),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47488),
            .ce(N__47851),
            .sr(N__46992));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_15_10_6  (
            .in0(N__48250),
            .in1(N__36429),
            .in2(_gnd_net_),
            .in3(N__36408),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47488),
            .ce(N__47851),
            .sr(N__46992));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_11_0  (
            .in0(N__41707),
            .in1(N__41678),
            .in2(_gnd_net_),
            .in3(N__48327),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_11_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_15_11_1  (
            .in0(N__48329),
            .in1(_gnd_net_),
            .in2(N__36765),
            .in3(N__41708),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47475),
            .ce(N__47862),
            .sr(N__47001));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_11_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_11_2  (
            .in0(N__36737),
            .in1(N__48328),
            .in2(_gnd_net_),
            .in3(N__36752),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(elapsed_time_ns_1_RNI4EOBB_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_11_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_15_11_3  (
            .in0(N__48331),
            .in1(_gnd_net_),
            .in2(N__36741),
            .in3(N__36738),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47475),
            .ce(N__47862),
            .sr(N__47001));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_11_4 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_11_4  (
            .in0(N__39164),
            .in1(N__36626),
            .in2(N__39189),
            .in3(N__36698),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_11_5 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_11_5  (
            .in0(N__36627),
            .in1(N__39165),
            .in2(N__36702),
            .in3(N__39185),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_11_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_11_6  (
            .in0(N__36661),
            .in1(N__48326),
            .in2(_gnd_net_),
            .in3(N__36677),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_15_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_15_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_15_11_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_15_11_7  (
            .in0(N__48330),
            .in1(_gnd_net_),
            .in2(N__36666),
            .in3(N__36662),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47475),
            .ce(N__47862),
            .sr(N__47001));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_12_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_12_3  (
            .in0(N__46148),
            .in1(N__46171),
            .in2(_gnd_net_),
            .in3(N__48325),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_15_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_15_12_4 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_15_12_4  (
            .in0(N__36983),
            .in1(N__46655),
            .in2(N__36966),
            .in3(N__36954),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_15_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_15_12_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36948),
            .in3(N__46558),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_15_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_15_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__46559),
            .in2(_gnd_net_),
            .in3(N__36935),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__39462),
            .in2(N__36920),
            .in3(N__36916),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__46230),
            .in2(_gnd_net_),
            .in3(N__36852),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__42507),
            .in2(_gnd_net_),
            .in3(N__36819),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__42519),
            .in2(_gnd_net_),
            .in3(N__36786),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__36783),
            .in2(_gnd_net_),
            .in3(N__36768),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__37203),
            .in2(_gnd_net_),
            .in3(N__37167),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__42543),
            .in2(_gnd_net_),
            .in3(N__37140),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(N__42531),
            .in2(_gnd_net_),
            .in3(N__37137),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__39300),
            .in2(_gnd_net_),
            .in3(N__37107),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__39321),
            .in2(_gnd_net_),
            .in3(N__37080),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__46335),
            .in2(_gnd_net_),
            .in3(N__37077),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__42144),
            .in2(_gnd_net_),
            .in3(N__37041),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__42153),
            .in2(_gnd_net_),
            .in3(N__36999),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__36996),
            .in2(_gnd_net_),
            .in3(N__36987),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__39639),
            .in2(_gnd_net_),
            .in3(N__37257),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__39621),
            .in2(_gnd_net_),
            .in3(N__37254),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__39306),
            .in2(_gnd_net_),
            .in3(N__37251),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__39612),
            .in2(_gnd_net_),
            .in3(N__37248),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__39312),
            .in2(_gnd_net_),
            .in3(N__37245),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__39327),
            .in2(_gnd_net_),
            .in3(N__37242),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__39645),
            .in2(_gnd_net_),
            .in3(N__37212),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__46188),
            .in2(_gnd_net_),
            .in3(N__37209),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__46287),
            .in2(_gnd_net_),
            .in3(N__37206),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__39630),
            .in2(_gnd_net_),
            .in3(N__37308),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__37506),
            .in2(_gnd_net_),
            .in3(N__37305),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__39516),
            .in2(_gnd_net_),
            .in3(N__37302),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__39507),
            .in2(_gnd_net_),
            .in3(N__37299),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__42135),
            .in2(_gnd_net_),
            .in3(N__37296),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__41316),
            .in2(_gnd_net_),
            .in3(N__37293),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37290),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_6 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_6  (
            .in0(N__40594),
            .in1(N__42932),
            .in2(N__37656),
            .in3(N__40175),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_16_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_16_7  (
            .in0(N__40174),
            .in1(N__40595),
            .in2(N__46323),
            .in3(N__37682),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_17_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_17_0  (
            .in0(N__42400),
            .in1(N__38012),
            .in2(_gnd_net_),
            .in3(N__37537),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43416),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_17_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_17_2  (
            .in0(N__42581),
            .in1(N__38014),
            .in2(_gnd_net_),
            .in3(N__37499),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_17_3 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_17_3  (
            .in0(N__38011),
            .in1(N__37471),
            .in2(_gnd_net_),
            .in3(N__39490),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_17_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_17_4  (
            .in0(N__46372),
            .in1(N__38013),
            .in2(_gnd_net_),
            .in3(N__37423),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_5  (
            .in0(N__40581),
            .in1(N__43391),
            .in2(N__40266),
            .in3(N__40291),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_17_6 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_17_6  (
            .in0(N__43132),
            .in1(N__37372),
            .in2(_gnd_net_),
            .in3(N__38015),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_17_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_17_7  (
            .in0(N__40228),
            .in1(N__40582),
            .in2(N__39452),
            .in3(N__39406),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_18_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_18_0  (
            .in0(N__40625),
            .in1(N__43473),
            .in2(N__40267),
            .in3(N__37917),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_18_1 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_18_1  (
            .in0(N__39365),
            .in1(N__46217),
            .in2(_gnd_net_),
            .in3(N__38039),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_18_2  (
            .in0(N__38034),
            .in1(N__43087),
            .in2(_gnd_net_),
            .in3(N__37775),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_18_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_18_3  (
            .in0(N__37742),
            .in1(N__38037),
            .in2(_gnd_net_),
            .in3(N__42959),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_18_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_18_4  (
            .in0(N__38035),
            .in1(N__43046),
            .in2(_gnd_net_),
            .in3(N__37712),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_18_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_18_5  (
            .in0(N__46318),
            .in1(N__37683),
            .in2(_gnd_net_),
            .in3(N__38040),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_18_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_18_6  (
            .in0(N__38038),
            .in1(N__42931),
            .in2(_gnd_net_),
            .in3(N__37655),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_18_7 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_18_7  (
            .in0(N__42997),
            .in1(N__37616),
            .in2(_gnd_net_),
            .in3(N__38036),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_19_0  (
            .in0(N__38017),
            .in1(N__42796),
            .in2(_gnd_net_),
            .in3(N__37574),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_1  (
            .in0(N__40611),
            .in1(N__46218),
            .in2(N__40268),
            .in3(N__39369),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_19_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_19_2  (
            .in0(N__43273),
            .in1(N__40610),
            .in2(_gnd_net_),
            .in3(N__38314),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_15_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_15_19_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_15_19_3  (
            .in0(N__40608),
            .in1(N__43346),
            .in2(_gnd_net_),
            .in3(N__38063),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_15_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_15_19_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_15_19_4  (
            .in0(N__38018),
            .in1(N__43471),
            .in2(_gnd_net_),
            .in3(N__37916),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_15_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_15_19_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_15_19_5  (
            .in0(N__40606),
            .in1(N__43426),
            .in2(_gnd_net_),
            .in3(N__37829),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_6  (
            .in0(N__43312),
            .in1(N__40609),
            .in2(_gnd_net_),
            .in3(N__37874),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_19_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_19_7  (
            .in0(N__40607),
            .in1(N__43390),
            .in2(_gnd_net_),
            .in3(N__40293),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_0 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_0  (
            .in0(N__40246),
            .in1(N__40565),
            .in2(N__37836),
            .in3(N__43427),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__40564),
            .in2(_gnd_net_),
            .in3(N__39411),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_20_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_20_7  (
            .in0(N__40566),
            .in1(N__40245),
            .in2(N__43280),
            .in3(N__38316),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_22_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__38248),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38226),
            .ce(),
            .sr(N__47063));
    defparam \delay_measurement_inst.start_timer_tr_LC_15_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_15_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_15_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38247),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38225),
            .ce(),
            .sr(N__47064));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_16_4_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_16_4_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_16_4_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_16_4_7  (
            .in0(_gnd_net_),
            .in1(N__38104),
            .in2(_gnd_net_),
            .in3(N__38212),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_16_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_16_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_16_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_16_5_2  (
            .in0(N__38390),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47550),
            .ce(),
            .sr(N__46957));
    defparam \phase_controller_inst2.stoper_tr.running_LC_16_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_16_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_16_5_3 .LUT_INIT=16'b1011000011111100;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_16_5_3  (
            .in0(N__38882),
            .in1(N__41283),
            .in2(N__38406),
            .in3(N__38366),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47550),
            .ce(),
            .sr(N__46957));
    defparam \phase_controller_inst2.start_timer_tr_LC_16_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_16_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_16_5_4 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_16_5_4  (
            .in0(N__38199),
            .in1(N__38187),
            .in2(N__38391),
            .in3(N__46467),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47550),
            .ce(),
            .sr(N__46957));
    defparam \phase_controller_inst2.state_2_LC_16_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_16_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_16_5_5 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_inst2.state_2_LC_16_5_5  (
            .in0(N__38173),
            .in1(N__38133),
            .in2(N__38457),
            .in3(N__39575),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47550),
            .ce(),
            .sr(N__46957));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_16_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_16_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_16_5_6 .LUT_INIT=16'b1111010100100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_16_5_6  (
            .in0(N__41282),
            .in1(N__38883),
            .in2(N__38367),
            .in3(N__38105),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47550),
            .ce(),
            .sr(N__46957));
    defparam \phase_controller_inst2.T12_LC_16_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.T12_LC_16_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T12_LC_16_5_7 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \phase_controller_inst2.T12_LC_16_5_7  (
            .in0(N__38455),
            .in1(N__38417),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47550),
            .ce(),
            .sr(N__46957));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_16_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_16_6_3 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_16_6_3  (
            .in0(N__38402),
            .in1(N__38361),
            .in2(_gnd_net_),
            .in3(N__38385),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_5  (
            .in0(_gnd_net_),
            .in1(N__41279),
            .in2(_gnd_net_),
            .in3(N__41258),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_16_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_16_6_6 .LUT_INIT=16'b1111110101011101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_16_6_6  (
            .in0(N__38360),
            .in1(N__41871),
            .in2(N__41853),
            .in3(N__38898),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_16_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_16_6_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_16_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38340),
            .in3(N__41280),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_7_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_7_0  (
            .in0(N__41495),
            .in1(N__41471),
            .in2(N__38328),
            .in3(N__38337),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_16_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_16_7_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_16_7_1  (
            .in0(N__38336),
            .in1(N__41496),
            .in2(N__41475),
            .in3(N__38324),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_2  (
            .in0(N__45279),
            .in1(N__45316),
            .in2(_gnd_net_),
            .in3(N__48228),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47535),
            .ce(N__46077),
            .sr(N__46966));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_16_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_16_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_16_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_16_7_3  (
            .in0(N__48225),
            .in1(N__44259),
            .in2(_gnd_net_),
            .in3(N__44298),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47535),
            .ce(N__46077),
            .sr(N__46966));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_16_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_16_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_16_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_16_7_4  (
            .in0(N__44617),
            .in1(N__44643),
            .in2(_gnd_net_),
            .in3(N__48229),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47535),
            .ce(N__46077),
            .sr(N__46966));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_16_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_16_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_16_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_16_7_5  (
            .in0(N__48226),
            .in1(N__44767),
            .in2(_gnd_net_),
            .in3(N__44205),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47535),
            .ce(N__46077),
            .sr(N__46966));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_16_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_16_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_16_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_16_7_6  (
            .in0(N__44805),
            .in1(N__44234),
            .in2(_gnd_net_),
            .in3(N__48230),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47535),
            .ce(N__46077),
            .sr(N__46966));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_16_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_16_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_16_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_16_7_7  (
            .in0(N__48227),
            .in1(N__45345),
            .in2(_gnd_net_),
            .in3(N__45370),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47535),
            .ce(N__46077),
            .sr(N__46966));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_16_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_16_8_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_16_8_0  (
            .in0(N__40715),
            .in1(N__38538),
            .in2(N__38532),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_16_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_16_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__38523),
            .in2(N__38514),
            .in3(N__40682),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_16_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_16_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__38505),
            .in2(N__38496),
            .in3(N__40658),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_16_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_16_8_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_16_8_3  (
            .in0(N__40643),
            .in1(N__38487),
            .in2(N__38481),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_16_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_16_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__38463),
            .in2(N__38472),
            .in3(N__41444),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_16_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_16_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__38637),
            .in2(N__38631),
            .in3(N__41430),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_16_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_16_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__38622),
            .in2(N__38616),
            .in3(N__41408),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_16_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_16_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__46095),
            .in2(N__38604),
            .in3(N__41393),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_16_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_16_9_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_16_9_0  (
            .in0(N__41379),
            .in1(N__38595),
            .in2(N__45027),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_16_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_16_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__44952),
            .in2(N__38589),
            .in3(N__41360),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_16_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_16_9_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_16_9_2  (
            .in0(N__41345),
            .in1(N__38580),
            .in2(N__38574),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_16_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_16_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__38565),
            .in2(N__38559),
            .in3(N__41330),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_16_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_16_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__46107),
            .in2(N__38550),
            .in3(N__41588),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_16_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_16_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_16_9_5  (
            .in0(N__41573),
            .in1(N__41667),
            .in2(N__38715),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_16_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_16_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_16_9_6  (
            .in0(N__41558),
            .in1(N__38697),
            .in2(N__38706),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_16_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_16_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__38691),
            .in2(N__38685),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_16_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_16_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__38676),
            .in2(N__38667),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_16_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_16_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__45255),
            .in2(N__45210),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_16_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_16_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__38652),
            .in2(N__38646),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_16_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_16_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__44940),
            .in2(N__44898),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_16_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_16_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__45504),
            .in2(N__45453),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_16_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_16_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__45441),
            .in2(N__45393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__41867),
            .in2(N__41733),
            .in3(N__38889),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38886),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_16_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_16_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__38868),
            .in2(N__38862),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_11_1  (
            .in0(N__47837),
            .in1(N__38822),
            .in2(_gnd_net_),
            .in3(N__38808),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__47489),
            .ce(),
            .sr(N__46993));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_16_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_16_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_16_11_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_16_11_2  (
            .in0(N__47841),
            .in1(N__38789),
            .in2(N__38805),
            .in3(N__38775),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__47489),
            .ce(),
            .sr(N__46993));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_16_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_16_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_16_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_16_11_3  (
            .in0(N__47838),
            .in1(N__38771),
            .in2(_gnd_net_),
            .in3(N__38757),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__47489),
            .ce(),
            .sr(N__46993));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_16_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_16_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_16_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_16_11_4  (
            .in0(N__47842),
            .in1(N__38753),
            .in2(_gnd_net_),
            .in3(N__38739),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__47489),
            .ce(),
            .sr(N__46993));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_16_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_16_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_16_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_16_11_5  (
            .in0(N__47839),
            .in1(N__38732),
            .in2(_gnd_net_),
            .in3(N__38718),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__47489),
            .ce(),
            .sr(N__46993));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_16_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_16_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_16_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_16_11_6  (
            .in0(N__47843),
            .in1(N__39041),
            .in2(_gnd_net_),
            .in3(N__39027),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__47489),
            .ce(),
            .sr(N__46993));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_16_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_16_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_16_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_16_11_7  (
            .in0(N__47840),
            .in1(N__39023),
            .in2(_gnd_net_),
            .in3(N__39009),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__47489),
            .ce(),
            .sr(N__46993));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_16_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_16_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_16_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_16_12_0  (
            .in0(N__47850),
            .in1(N__39005),
            .in2(_gnd_net_),
            .in3(N__38991),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__47476),
            .ce(),
            .sr(N__47002));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_16_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_16_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_16_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_16_12_1  (
            .in0(N__47777),
            .in1(N__38987),
            .in2(_gnd_net_),
            .in3(N__38973),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__47476),
            .ce(),
            .sr(N__47002));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_16_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_16_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_16_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_16_12_2  (
            .in0(N__47847),
            .in1(N__38969),
            .in2(_gnd_net_),
            .in3(N__38955),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__47476),
            .ce(),
            .sr(N__47002));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_16_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_16_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_16_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_16_12_3  (
            .in0(N__47778),
            .in1(N__38951),
            .in2(_gnd_net_),
            .in3(N__38937),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__47476),
            .ce(),
            .sr(N__47002));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_16_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_16_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_16_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_16_12_4  (
            .in0(N__47848),
            .in1(N__38933),
            .in2(_gnd_net_),
            .in3(N__38919),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__47476),
            .ce(),
            .sr(N__47002));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_16_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_16_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_16_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_16_12_5  (
            .in0(N__47779),
            .in1(N__38915),
            .in2(_gnd_net_),
            .in3(N__38901),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__47476),
            .ce(),
            .sr(N__47002));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_16_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_16_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_16_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_16_12_6  (
            .in0(N__47849),
            .in1(N__39206),
            .in2(_gnd_net_),
            .in3(N__39192),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__47476),
            .ce(),
            .sr(N__47002));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_12_7  (
            .in0(N__47780),
            .in1(N__39184),
            .in2(_gnd_net_),
            .in3(N__39168),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__47476),
            .ce(),
            .sr(N__47002));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_16_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_16_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_16_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_16_13_0  (
            .in0(N__47833),
            .in1(N__39163),
            .in2(_gnd_net_),
            .in3(N__39147),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__47464),
            .ce(),
            .sr(N__47008));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_16_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_16_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_16_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_16_13_1  (
            .in0(N__47819),
            .in1(N__42231),
            .in2(_gnd_net_),
            .in3(N__39144),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__47464),
            .ce(),
            .sr(N__47008));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_16_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_16_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_16_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_16_13_2  (
            .in0(N__47834),
            .in1(N__42192),
            .in2(_gnd_net_),
            .in3(N__39141),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__47464),
            .ce(),
            .sr(N__47008));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_16_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_16_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_16_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_16_13_3  (
            .in0(N__47820),
            .in1(N__39133),
            .in2(_gnd_net_),
            .in3(N__39117),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__47464),
            .ce(),
            .sr(N__47008));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_16_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_16_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_16_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_16_13_4  (
            .in0(N__47835),
            .in1(N__39112),
            .in2(_gnd_net_),
            .in3(N__39096),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__47464),
            .ce(),
            .sr(N__47008));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_16_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_16_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_16_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_16_13_5  (
            .in0(N__47821),
            .in1(N__39083),
            .in2(_gnd_net_),
            .in3(N__39069),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__47464),
            .ce(),
            .sr(N__47008));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_16_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_16_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_16_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_16_13_6  (
            .in0(N__47836),
            .in1(N__39059),
            .in2(_gnd_net_),
            .in3(N__39045),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__47464),
            .ce(),
            .sr(N__47008));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_16_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_16_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_16_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_16_13_7  (
            .in0(N__47822),
            .in1(N__45854),
            .in2(_gnd_net_),
            .in3(N__39291),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__47464),
            .ce(),
            .sr(N__47008));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_16_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_16_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_16_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_16_14_0  (
            .in0(N__47829),
            .in1(N__45839),
            .in2(_gnd_net_),
            .in3(N__39288),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__47456),
            .ce(),
            .sr(N__47014));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_16_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_16_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_16_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_16_14_1  (
            .in0(N__47826),
            .in1(N__45926),
            .in2(_gnd_net_),
            .in3(N__39285),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__47456),
            .ce(),
            .sr(N__47014));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_16_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_16_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_16_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_16_14_2  (
            .in0(N__47830),
            .in1(N__45953),
            .in2(_gnd_net_),
            .in3(N__39282),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__47456),
            .ce(),
            .sr(N__47014));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_16_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_16_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_16_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_16_14_3  (
            .in0(N__47827),
            .in1(N__46037),
            .in2(_gnd_net_),
            .in3(N__39279),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__47456),
            .ce(),
            .sr(N__47014));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_16_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_16_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_16_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_16_14_4  (
            .in0(N__47831),
            .in1(N__46013),
            .in2(_gnd_net_),
            .in3(N__39276),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__47456),
            .ce(),
            .sr(N__47014));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_16_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_16_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_16_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_16_14_5  (
            .in0(N__47828),
            .in1(N__39257),
            .in2(_gnd_net_),
            .in3(N__39243),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__47456),
            .ce(),
            .sr(N__47014));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_16_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_16_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_16_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_16_14_6  (
            .in0(N__47832),
            .in1(N__39224),
            .in2(_gnd_net_),
            .in3(N__39240),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47456),
            .ce(),
            .sr(N__47014));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43710),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__43231),
            .sr(N__47021));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39480),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_16_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_16_15_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_16_15_7  (
            .in0(N__39453),
            .in1(N__40629),
            .in2(N__40271),
            .in3(N__39407),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_16_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_16_16_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_16_16_0  (
            .in0(N__40596),
            .in1(N__46210),
            .in2(N__40269),
            .in3(N__39364),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42913),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42694),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42947),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43029),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42732),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_16_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_16_6  (
            .in0(N__40597),
            .in1(N__40292),
            .in2(N__40270),
            .in3(N__43392),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42874),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43114),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43452),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43069),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42980),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.T01_LC_16_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.T01_LC_16_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T01_LC_16_17_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst2.T01_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__39527),
            .in2(_gnd_net_),
            .in3(N__39599),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47435),
            .ce(),
            .sr(N__47033));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43372),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43334),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43254),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_21_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__41307),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_17_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_17_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_17_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_17_5_3  (
            .in0(N__44251),
            .in1(N__44297),
            .in2(_gnd_net_),
            .in3(N__48189),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47554),
            .ce(N__47824),
            .sr(N__46955));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_17_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_17_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_17_6_0 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_17_6_0  (
            .in0(N__41281),
            .in1(N__41259),
            .in2(N__40716),
            .in3(N__42122),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47551),
            .ce(),
            .sr(N__46958));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_17_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_17_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_17_6_5  (
            .in0(N__40738),
            .in1(N__41247),
            .in2(_gnd_net_),
            .in3(N__41186),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(N__40711),
            .in2(N__40692),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_7_1  (
            .in0(N__42092),
            .in1(N__40683),
            .in2(_gnd_net_),
            .in3(N__40671),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__47545),
            .ce(),
            .sr(N__46961));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_7_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_7_2  (
            .in0(N__42096),
            .in1(N__40668),
            .in2(N__40662),
            .in3(N__40647),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__47545),
            .ce(),
            .sr(N__46961));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_7_3  (
            .in0(N__42093),
            .in1(N__40644),
            .in2(_gnd_net_),
            .in3(N__40632),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__47545),
            .ce(),
            .sr(N__46961));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_7_4  (
            .in0(N__42097),
            .in1(N__41445),
            .in2(_gnd_net_),
            .in3(N__41433),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__47545),
            .ce(),
            .sr(N__46961));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_7_5  (
            .in0(N__42094),
            .in1(N__41426),
            .in2(_gnd_net_),
            .in3(N__41412),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__47545),
            .ce(),
            .sr(N__46961));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_7_6  (
            .in0(N__42098),
            .in1(N__41409),
            .in2(_gnd_net_),
            .in3(N__41397),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__47545),
            .ce(),
            .sr(N__46961));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_7_7  (
            .in0(N__42095),
            .in1(N__41394),
            .in2(_gnd_net_),
            .in3(N__41382),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__47545),
            .ce(),
            .sr(N__46961));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_8_0  (
            .in0(N__42106),
            .in1(N__41378),
            .in2(_gnd_net_),
            .in3(N__41364),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__47536),
            .ce(),
            .sr(N__46967));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_8_1  (
            .in0(N__42099),
            .in1(N__41361),
            .in2(_gnd_net_),
            .in3(N__41349),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__47536),
            .ce(),
            .sr(N__46967));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_8_2  (
            .in0(N__42103),
            .in1(N__41346),
            .in2(_gnd_net_),
            .in3(N__41334),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__47536),
            .ce(),
            .sr(N__46967));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_8_3  (
            .in0(N__42100),
            .in1(N__41331),
            .in2(_gnd_net_),
            .in3(N__41319),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__47536),
            .ce(),
            .sr(N__46967));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_8_4  (
            .in0(N__42104),
            .in1(N__41589),
            .in2(_gnd_net_),
            .in3(N__41577),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__47536),
            .ce(),
            .sr(N__46967));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_8_5  (
            .in0(N__42101),
            .in1(N__41574),
            .in2(_gnd_net_),
            .in3(N__41562),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__47536),
            .ce(),
            .sr(N__46967));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_8_6  (
            .in0(N__42105),
            .in1(N__41559),
            .in2(_gnd_net_),
            .in3(N__41547),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__47536),
            .ce(),
            .sr(N__46967));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_8_7  (
            .in0(N__42102),
            .in1(N__41542),
            .in2(_gnd_net_),
            .in3(N__41526),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__47536),
            .ce(),
            .sr(N__46967));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_9_0  (
            .in0(N__42107),
            .in1(N__41513),
            .in2(_gnd_net_),
            .in3(N__41499),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__47526),
            .ce(),
            .sr(N__46973));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_9_1  (
            .in0(N__42111),
            .in1(N__41494),
            .in2(_gnd_net_),
            .in3(N__41478),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__47526),
            .ce(),
            .sr(N__46973));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_9_2  (
            .in0(N__42108),
            .in1(N__41470),
            .in2(_gnd_net_),
            .in3(N__41454),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__47526),
            .ce(),
            .sr(N__46973));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_17_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_17_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_17_9_3  (
            .in0(N__42112),
            .in1(N__45227),
            .in2(_gnd_net_),
            .in3(N__41451),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__47526),
            .ce(),
            .sr(N__46973));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_17_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_17_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_17_9_4  (
            .in0(N__42109),
            .in1(N__45243),
            .in2(_gnd_net_),
            .in3(N__41448),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__47526),
            .ce(),
            .sr(N__46973));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_17_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_17_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_17_9_5  (
            .in0(N__42113),
            .in1(N__41656),
            .in2(_gnd_net_),
            .in3(N__41640),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__47526),
            .ce(),
            .sr(N__46973));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_17_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_17_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_17_9_6  (
            .in0(N__42110),
            .in1(N__41632),
            .in2(_gnd_net_),
            .in3(N__41613),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__47526),
            .ce(),
            .sr(N__46973));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_17_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_17_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_17_9_7  (
            .in0(N__42114),
            .in1(N__44915),
            .in2(_gnd_net_),
            .in3(N__41610),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__47526),
            .ce(),
            .sr(N__46973));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_17_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_17_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_17_10_0  (
            .in0(N__42115),
            .in1(N__44931),
            .in2(_gnd_net_),
            .in3(N__41607),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__47515),
            .ce(),
            .sr(N__46980));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_17_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_17_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_17_10_1  (
            .in0(N__42119),
            .in1(N__45479),
            .in2(_gnd_net_),
            .in3(N__41604),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__47515),
            .ce(),
            .sr(N__46980));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_17_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_17_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_17_10_2  (
            .in0(N__42116),
            .in1(N__45495),
            .in2(_gnd_net_),
            .in3(N__41601),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__47515),
            .ce(),
            .sr(N__46980));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_17_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_17_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_17_10_3  (
            .in0(N__42120),
            .in1(N__45428),
            .in2(_gnd_net_),
            .in3(N__41598),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__47515),
            .ce(),
            .sr(N__46980));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_17_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_17_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_17_10_4  (
            .in0(N__42117),
            .in1(N__45410),
            .in2(_gnd_net_),
            .in3(N__41595),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__47515),
            .ce(),
            .sr(N__46980));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_17_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_17_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_17_10_5  (
            .in0(N__42121),
            .in1(N__41755),
            .in2(_gnd_net_),
            .in3(N__41592),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__47515),
            .ce(),
            .sr(N__46980));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_17_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_17_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_17_10_6  (
            .in0(N__42118),
            .in1(N__41775),
            .in2(_gnd_net_),
            .in3(N__41958),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47515),
            .ce(),
            .sr(N__46980));
    defparam \phase_controller_inst2.T23_LC_17_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.T23_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T23_LC_17_10_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst2.T23_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__41882),
            .in2(_gnd_net_),
            .in3(N__41944),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47515),
            .ce(),
            .sr(N__46980));
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_17_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_17_11_0 .LUT_INIT=16'b0010101100001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_17_11_0  (
            .in0(N__41772),
            .in1(N__41748),
            .in2(N__41724),
            .in3(N__41786),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_17_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_17_11_1 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_17_11_1  (
            .in0(N__41785),
            .in1(N__41773),
            .in2(N__41756),
            .in3(N__41719),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_17_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_17_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_30_LC_17_11_2  (
            .in0(N__48340),
            .in1(N__41838),
            .in2(_gnd_net_),
            .in3(N__41805),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47501),
            .ce(N__46080),
            .sr(N__46986));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_17_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_17_11_3 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_17_11_3  (
            .in0(N__41787),
            .in1(N__41774),
            .in2(N__41757),
            .in3(N__41723),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_17_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_17_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_31_LC_17_11_6  (
            .in0(N__48341),
            .in1(N__44716),
            .in2(_gnd_net_),
            .in3(N__44325),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47501),
            .ce(N__46080),
            .sr(N__46986));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_17_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_17_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_17_11_7  (
            .in0(N__41709),
            .in1(N__41682),
            .in2(_gnd_net_),
            .in3(N__48342),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47501),
            .ce(N__46080),
            .sr(N__46986));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_12_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_12_1  (
            .in0(N__42242),
            .in1(N__42190),
            .in2(N__42212),
            .in3(N__42229),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_12_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_12_5  (
            .in0(N__42284),
            .in1(N__48294),
            .in2(_gnd_net_),
            .in3(N__42296),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(elapsed_time_ns_1_RNI2COBB_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_17_12_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_17_12_6  (
            .in0(N__48295),
            .in1(N__42285),
            .in2(N__42255),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47490),
            .ce(N__47815),
            .sr(N__46994));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_17_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_17_12_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_17_12_7  (
            .in0(N__45318),
            .in1(N__45271),
            .in2(_gnd_net_),
            .in3(N__48296),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47490),
            .ce(N__47815),
            .sr(N__46994));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_13_0 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_13_0  (
            .in0(N__42243),
            .in1(N__42230),
            .in2(N__42213),
            .in3(N__42191),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_13_6 .LUT_INIT=16'b1011001010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_13_6  (
            .in0(N__45905),
            .in1(N__45949),
            .in2(N__45978),
            .in3(N__45925),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42604),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42651),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_14_3  (
            .in0(N__43303),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42820),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42777),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42427),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42472),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_17_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_17_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_17_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__43166),
            .in2(N__43679),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47457),
            .ce(N__43233),
            .sr(N__47015));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_17_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_17_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_17_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__43706),
            .in2(N__43650),
            .in3(N__42456),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47457),
            .ce(N__43233),
            .sr(N__47015));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_17_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_17_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_17_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__43680),
            .in2(N__43619),
            .in3(N__42411),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47457),
            .ce(N__43233),
            .sr(N__47015));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_17_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_17_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_17_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__43649),
            .in2(N__43589),
            .in3(N__42363),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47457),
            .ce(N__43233),
            .sr(N__47015));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_17_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_17_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_17_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__43559),
            .in2(N__43620),
            .in3(N__42321),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47457),
            .ce(N__43233),
            .sr(N__47015));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_17_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_17_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_17_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__43532),
            .in2(N__43590),
            .in3(N__42804),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47457),
            .ce(N__43233),
            .sr(N__47015));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_17_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_17_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_17_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__43560),
            .in2(N__43505),
            .in3(N__42759),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47457),
            .ce(N__43233),
            .sr(N__47015));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_17_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_17_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_17_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__43955),
            .in2(N__43536),
            .in3(N__42717),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47457),
            .ce(N__43233),
            .sr(N__47015));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_17_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_17_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_17_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__43928),
            .in2(N__43506),
            .in3(N__42678),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47447),
            .ce(N__43232),
            .sr(N__47022));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_17_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_17_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_17_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__43907),
            .in2(N__43962),
            .in3(N__42675),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47447),
            .ce(N__43232),
            .sr(N__47022));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_17_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_17_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_17_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__43929),
            .in2(N__43884),
            .in3(N__42624),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47447),
            .ce(N__43232),
            .sr(N__47022));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_17_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_17_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_17_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__43908),
            .in2(N__43856),
            .in3(N__42585),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47447),
            .ce(N__43232),
            .sr(N__47022));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_17_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_17_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_17_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__43883),
            .in2(N__43826),
            .in3(N__42546),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47447),
            .ce(N__43232),
            .sr(N__47022));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_17_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_17_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_17_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__43796),
            .in2(N__43857),
            .in3(N__43098),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47447),
            .ce(N__43232),
            .sr(N__47022));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_17_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_17_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_17_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__43769),
            .in2(N__43827),
            .in3(N__43053),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47447),
            .ce(N__43232),
            .sr(N__47022));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_17_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_17_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_17_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__43797),
            .in2(N__43743),
            .in3(N__43011),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47447),
            .ce(N__43232),
            .sr(N__47022));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_17_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_17_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_17_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__44174),
            .in2(N__43773),
            .in3(N__42969),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47441),
            .ce(N__43230),
            .sr(N__47028));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_17_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_17_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_17_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__43742),
            .in2(N__44147),
            .in3(N__42936),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47441),
            .ce(N__43230),
            .sr(N__47028));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_17_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_17_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_17_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__44120),
            .in2(N__44178),
            .in3(N__42897),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47441),
            .ce(N__43230),
            .sr(N__47028));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_17_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_17_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_17_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__44096),
            .in2(N__44148),
            .in3(N__42861),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47441),
            .ce(N__43230),
            .sr(N__47028));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_17_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_17_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_17_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__44121),
            .in2(N__44072),
            .in3(N__42858),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47441),
            .ce(N__43230),
            .sr(N__47028));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_17_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_17_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_17_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__44045),
            .in2(N__44100),
            .in3(N__42855),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47441),
            .ce(N__43230),
            .sr(N__47028));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_17_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_17_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_17_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__44021),
            .in2(N__44073),
            .in3(N__43431),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47441),
            .ce(N__43230),
            .sr(N__47028));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_17_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_17_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_17_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__44046),
            .in2(N__43994),
            .in3(N__43395),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47441),
            .ce(N__43230),
            .sr(N__47028));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_17_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_17_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__44570),
            .in2(N__44025),
            .in3(N__43356),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47436),
            .ce(N__43228),
            .sr(N__47034));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_17_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_17_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__43995),
            .in2(N__44543),
            .in3(N__43323),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47436),
            .ce(N__43228),
            .sr(N__47034));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_17_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_17_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__44517),
            .in2(N__44574),
            .in3(N__43284),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47436),
            .ce(N__43228),
            .sr(N__47034));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_17_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_17_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__44379),
            .in2(N__44544),
            .in3(N__43236),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47436),
            .ce(N__43228),
            .sr(N__47034));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_17_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_17_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43203),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_17_19_0  (
            .in0(N__44489),
            .in1(N__43162),
            .in2(_gnd_net_),
            .in3(N__43143),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__47432),
            .ce(N__44356),
            .sr(N__47040));
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_17_19_1  (
            .in0(N__44485),
            .in1(N__43702),
            .in2(_gnd_net_),
            .in3(N__43683),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__47432),
            .ce(N__44356),
            .sr(N__47040));
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_17_19_2  (
            .in0(N__44490),
            .in1(N__43672),
            .in2(_gnd_net_),
            .in3(N__43653),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__47432),
            .ce(N__44356),
            .sr(N__47040));
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_17_19_3  (
            .in0(N__44486),
            .in1(N__43639),
            .in2(_gnd_net_),
            .in3(N__43623),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__47432),
            .ce(N__44356),
            .sr(N__47040));
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_17_19_4  (
            .in0(N__44491),
            .in1(N__43607),
            .in2(_gnd_net_),
            .in3(N__43593),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__47432),
            .ce(N__44356),
            .sr(N__47040));
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_17_19_5  (
            .in0(N__44487),
            .in1(N__43577),
            .in2(_gnd_net_),
            .in3(N__43563),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__47432),
            .ce(N__44356),
            .sr(N__47040));
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_17_19_6  (
            .in0(N__44492),
            .in1(N__43553),
            .in2(_gnd_net_),
            .in3(N__43539),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__47432),
            .ce(N__44356),
            .sr(N__47040));
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_17_19_7  (
            .in0(N__44488),
            .in1(N__43525),
            .in2(_gnd_net_),
            .in3(N__43509),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__47432),
            .ce(N__44356),
            .sr(N__47040));
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_17_20_0  (
            .in0(N__44496),
            .in1(N__43492),
            .in2(_gnd_net_),
            .in3(N__43476),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__47428),
            .ce(N__44363),
            .sr(N__47045));
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_17_20_1  (
            .in0(N__44477),
            .in1(N__43954),
            .in2(_gnd_net_),
            .in3(N__43932),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__47428),
            .ce(N__44363),
            .sr(N__47045));
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_17_20_2  (
            .in0(N__44493),
            .in1(N__43927),
            .in2(_gnd_net_),
            .in3(N__43911),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__47428),
            .ce(N__44363),
            .sr(N__47045));
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_17_20_3  (
            .in0(N__44474),
            .in1(N__43901),
            .in2(_gnd_net_),
            .in3(N__43887),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__47428),
            .ce(N__44363),
            .sr(N__47045));
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_17_20_4  (
            .in0(N__44494),
            .in1(N__43879),
            .in2(_gnd_net_),
            .in3(N__43860),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__47428),
            .ce(N__44363),
            .sr(N__47045));
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_17_20_5  (
            .in0(N__44475),
            .in1(N__43844),
            .in2(_gnd_net_),
            .in3(N__43830),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__47428),
            .ce(N__44363),
            .sr(N__47045));
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_17_20_6  (
            .in0(N__44495),
            .in1(N__43814),
            .in2(_gnd_net_),
            .in3(N__43800),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__47428),
            .ce(N__44363),
            .sr(N__47045));
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_17_20_7  (
            .in0(N__44476),
            .in1(N__43790),
            .in2(_gnd_net_),
            .in3(N__43776),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__47428),
            .ce(N__44363),
            .sr(N__47045));
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_17_21_0  (
            .in0(N__44470),
            .in1(N__43762),
            .in2(_gnd_net_),
            .in3(N__43746),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__47427),
            .ce(N__44355),
            .sr(N__47051));
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_17_21_1  (
            .in0(N__44481),
            .in1(N__43732),
            .in2(_gnd_net_),
            .in3(N__43713),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__47427),
            .ce(N__44355),
            .sr(N__47051));
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_17_21_2  (
            .in0(N__44471),
            .in1(N__44167),
            .in2(_gnd_net_),
            .in3(N__44151),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__47427),
            .ce(N__44355),
            .sr(N__47051));
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_17_21_3  (
            .in0(N__44482),
            .in1(N__44140),
            .in2(_gnd_net_),
            .in3(N__44124),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__47427),
            .ce(N__44355),
            .sr(N__47051));
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_17_21_4  (
            .in0(N__44472),
            .in1(N__44119),
            .in2(_gnd_net_),
            .in3(N__44103),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__47427),
            .ce(N__44355),
            .sr(N__47051));
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_17_21_5  (
            .in0(N__44483),
            .in1(N__44095),
            .in2(_gnd_net_),
            .in3(N__44076),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__47427),
            .ce(N__44355),
            .sr(N__47051));
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_17_21_6  (
            .in0(N__44473),
            .in1(N__44065),
            .in2(_gnd_net_),
            .in3(N__44049),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__47427),
            .ce(N__44355),
            .sr(N__47051));
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_17_21_7  (
            .in0(N__44484),
            .in1(N__44044),
            .in2(_gnd_net_),
            .in3(N__44028),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__47427),
            .ce(N__44355),
            .sr(N__47051));
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_17_22_0  (
            .in0(N__44497),
            .in1(N__44014),
            .in2(_gnd_net_),
            .in3(N__43998),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__47426),
            .ce(N__44364),
            .sr(N__47055));
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_17_22_1  (
            .in0(N__44478),
            .in1(N__43987),
            .in2(_gnd_net_),
            .in3(N__43965),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__47426),
            .ce(N__44364),
            .sr(N__47055));
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_17_22_2  (
            .in0(N__44498),
            .in1(N__44563),
            .in2(_gnd_net_),
            .in3(N__44547),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__47426),
            .ce(N__44364),
            .sr(N__47055));
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_17_22_3  (
            .in0(N__44479),
            .in1(N__44536),
            .in2(_gnd_net_),
            .in3(N__44520),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__47426),
            .ce(N__44364),
            .sr(N__47055));
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_17_22_4  (
            .in0(N__44499),
            .in1(N__44516),
            .in2(_gnd_net_),
            .in3(N__44502),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__47426),
            .ce(N__44364),
            .sr(N__47055));
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_17_22_5  (
            .in0(N__44480),
            .in1(N__44378),
            .in2(_gnd_net_),
            .in3(N__44382),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47426),
            .ce(N__44364),
            .sr(N__47055));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_5_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_5_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_5_4  (
            .in0(N__44320),
            .in1(N__44721),
            .in2(_gnd_net_),
            .in3(N__48188),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_5_5  (
            .in0(N__48187),
            .in1(N__44255),
            .in2(_gnd_net_),
            .in3(N__44296),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_18_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_18_6_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_18_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_18_6_0  (
            .in0(N__48042),
            .in1(N__44808),
            .in2(_gnd_net_),
            .in3(N__44233),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_18_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_18_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_18_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_18_6_1  (
            .in0(N__44200),
            .in1(N__44769),
            .in2(_gnd_net_),
            .in3(N__48043),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_18_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_18_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_18_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_18_6_6  (
            .in0(N__48041),
            .in1(N__45010),
            .in2(_gnd_net_),
            .in3(N__44990),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_18_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_18_7_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_18_7_0  (
            .in0(_gnd_net_),
            .in1(N__48448),
            .in2(_gnd_net_),
            .in3(N__45369),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_18_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_18_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_18_7_2  (
            .in0(N__44886),
            .in1(N__44976),
            .in2(N__44847),
            .in3(N__45051),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_18_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_18_7_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_18_7_3  (
            .in0(N__44806),
            .in1(N__44754),
            .in2(N__44730),
            .in3(N__44727),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_4 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_4  (
            .in0(N__44717),
            .in1(N__44676),
            .in2(N__44664),
            .in3(N__44649),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_5  (
            .in0(N__45052),
            .in1(_gnd_net_),
            .in2(N__44661),
            .in3(N__45079),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_18_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_18_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_18_7_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_18_7_6  (
            .in0(N__45586),
            .in1(N__45648),
            .in2(_gnd_net_),
            .in3(N__44658),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_7_7  (
            .in0(N__44642),
            .in1(N__44616),
            .in2(_gnd_net_),
            .in3(N__48044),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_18_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_18_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_18_8_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_26_LC_18_8_1  (
            .in0(N__45543),
            .in1(N__48073),
            .in2(_gnd_net_),
            .in3(N__45561),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47546),
            .ce(N__47873),
            .sr(N__46962));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_18_8_5  (
            .in0(N__44638),
            .in1(N__44622),
            .in2(_gnd_net_),
            .in3(N__48074),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47546),
            .ce(N__47873),
            .sr(N__46962));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_18_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_18_9_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_18_9_0  (
            .in0(N__45242),
            .in1(N__45223),
            .in2(N__45096),
            .in3(N__45147),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_1  (
            .in0(N__45146),
            .in1(N__45241),
            .in2(N__45228),
            .in3(N__45092),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_18_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_18_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_18_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_20_LC_18_9_2  (
            .in0(N__48184),
            .in1(N__45193),
            .in2(_gnd_net_),
            .in3(N__45165),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47537),
            .ce(N__46079),
            .sr(N__46968));
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_18_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_18_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_18_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_21_LC_18_9_5  (
            .in0(N__45138),
            .in1(N__48186),
            .in2(_gnd_net_),
            .in3(N__45117),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47537),
            .ce(N__46079),
            .sr(N__46968));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_18_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_18_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_18_9_6  (
            .in0(N__48185),
            .in1(N__45080),
            .in2(_gnd_net_),
            .in3(N__45060),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47537),
            .ce(N__46079),
            .sr(N__46968));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_18_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_18_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_18_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_18_9_7  (
            .in0(N__45011),
            .in1(N__44991),
            .in2(_gnd_net_),
            .in3(N__48120),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47537),
            .ce(N__46079),
            .sr(N__46968));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_10_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_10_0  (
            .in0(N__44930),
            .in1(N__45677),
            .in2(N__44916),
            .in3(N__45708),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_18_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_18_10_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_18_10_1  (
            .in0(N__45707),
            .in1(N__44929),
            .in2(N__45681),
            .in3(N__44914),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_18_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_18_10_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_18_10_2  (
            .in0(N__45541),
            .in1(N__48118),
            .in2(_gnd_net_),
            .in3(N__45557),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_18_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_18_10_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_26_LC_18_10_3  (
            .in0(N__48119),
            .in1(_gnd_net_),
            .in2(N__45546),
            .in3(N__45542),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47527),
            .ce(N__46081),
            .sr(N__46974));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_18_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_18_10_4 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_18_10_4  (
            .in0(N__45461),
            .in1(N__45478),
            .in2(N__45696),
            .in3(N__45493),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_10_5 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_10_5  (
            .in0(N__45494),
            .in1(N__45692),
            .in2(N__45480),
            .in3(N__45462),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_11_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_11_0  (
            .in0(N__45717),
            .in1(N__45726),
            .in2(N__45429),
            .in3(N__45409),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_18_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_18_11_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_18_11_1  (
            .in0(N__45725),
            .in1(N__45427),
            .in2(N__45411),
            .in3(N__45716),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_18_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_18_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_18_11_3  (
            .in0(N__48257),
            .in1(N__45344),
            .in2(_gnd_net_),
            .in3(N__45377),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_11_4  (
            .in0(N__45275),
            .in1(N__45317),
            .in2(_gnd_net_),
            .in3(N__48256),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_18_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_18_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_18_12_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_28_LC_18_12_0  (
            .in0(N__45597),
            .in1(N__48301),
            .in2(_gnd_net_),
            .in3(N__45612),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47502),
            .ce(N__46083),
            .sr(N__46987));
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_18_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_18_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_18_12_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_29_LC_18_12_1  (
            .in0(N__48298),
            .in1(N__48405),
            .in2(_gnd_net_),
            .in3(N__48377),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47502),
            .ce(N__46083),
            .sr(N__46987));
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_18_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_18_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_18_12_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_24_LC_18_12_2  (
            .in0(N__46509),
            .in1(N__48299),
            .in2(_gnd_net_),
            .in3(N__45741),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47502),
            .ce(N__46083),
            .sr(N__46987));
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_18_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_18_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_27_LC_18_12_3  (
            .in0(N__48297),
            .in1(N__45666),
            .in2(_gnd_net_),
            .in3(N__45651),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47502),
            .ce(N__46083),
            .sr(N__46987));
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_18_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_18_12_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_25_LC_18_12_6  (
            .in0(N__45786),
            .in1(N__48300),
            .in2(_gnd_net_),
            .in3(N__45804),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47502),
            .ce(N__46083),
            .sr(N__46987));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_18_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_18_13_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_18_13_0  (
            .in0(N__45649),
            .in1(N__48258),
            .in2(_gnd_net_),
            .in3(N__45665),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_18_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_18_13_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_27_LC_18_13_1  (
            .in0(N__48260),
            .in1(_gnd_net_),
            .in2(N__45654),
            .in3(N__45650),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47491),
            .ce(N__47811),
            .sr(N__46995));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_13_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_13_2  (
            .in0(N__45595),
            .in1(N__48259),
            .in2(_gnd_net_),
            .in3(N__45611),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_18_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_18_13_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_28_LC_18_13_3  (
            .in0(N__48261),
            .in1(_gnd_net_),
            .in2(N__45600),
            .in3(N__45596),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47491),
            .ce(N__47811),
            .sr(N__46995));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_18_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_18_13_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_18_13_4  (
            .in0(N__45998),
            .in1(N__46044),
            .in2(N__46023),
            .in3(N__47891),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_13_5 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_13_5  (
            .in0(N__46043),
            .in1(N__46022),
            .in2(N__47895),
            .in3(N__45999),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_13_7 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_13_7  (
            .in0(N__45977),
            .in1(N__45957),
            .in2(N__45933),
            .in3(N__45906),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_14_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_14_0  (
            .in0(N__45750),
            .in1(N__46476),
            .in2(N__45864),
            .in3(N__45835),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_14_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_14_1  (
            .in0(N__46475),
            .in1(N__45863),
            .in2(N__45840),
            .in3(N__45749),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_18_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_18_14_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_18_14_2  (
            .in0(N__45781),
            .in1(N__48253),
            .in2(_gnd_net_),
            .in3(N__45800),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_18_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_18_14_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_25_LC_18_14_3  (
            .in0(N__48255),
            .in1(_gnd_net_),
            .in2(N__45789),
            .in3(N__45782),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47477),
            .ce(N__47823),
            .sr(N__47003));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_18_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_18_14_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_18_14_4  (
            .in0(N__46501),
            .in1(N__48252),
            .in2(_gnd_net_),
            .in3(N__45737),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(elapsed_time_ns_1_RNI2DPBB_0_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_18_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_18_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_18_14_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_24_LC_18_14_5  (
            .in0(N__48254),
            .in1(_gnd_net_),
            .in2(N__46512),
            .in3(N__46502),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47477),
            .ce(N__47823),
            .sr(N__47003));
    defparam \phase_controller_inst1.start_timer_tr_LC_18_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_18_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_18_15_2 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_18_15_2  (
            .in0(N__46455),
            .in1(N__46413),
            .in2(N__46592),
            .in3(N__46398),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47465),
            .ce(),
            .sr(N__47009));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_18_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_18_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_18_15_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_18_15_6  (
            .in0(N__46587),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47465),
            .ce(),
            .sr(N__47009));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46353),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46300),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46248),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46204),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_20_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_20_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_20_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_20_8_1  (
            .in0(N__46176),
            .in1(N__46152),
            .in2(_gnd_net_),
            .in3(N__48305),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47555),
            .ce(N__46082),
            .sr(N__46963));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_20_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_20_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_20_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_20_8_7  (
            .in0(N__48421),
            .in1(N__48465),
            .in2(_gnd_net_),
            .in3(N__48306),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47555),
            .ce(N__46082),
            .sr(N__46963));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_20_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_20_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_20_9_4  (
            .in0(N__48425),
            .in1(N__48464),
            .in2(_gnd_net_),
            .in3(N__48293),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_20_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_20_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_20_10_3  (
            .in0(N__48400),
            .in1(N__48376),
            .in2(_gnd_net_),
            .in3(N__48262),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_6  (
            .in0(N__48401),
            .in1(N__48378),
            .in2(_gnd_net_),
            .in3(N__48338),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47528),
            .ce(N__47735),
            .sr(N__46988));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_4  (
            .in0(_gnd_net_),
            .in1(N__46650),
            .in2(_gnd_net_),
            .in3(N__46593),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_LC_20_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_20_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_20_14_4 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_20_14_4  (
            .in0(N__46651),
            .in1(N__47583),
            .in2(N__46608),
            .in3(N__46536),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47503),
            .ce(),
            .sr(N__47004));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5  (
            .in0(N__46637),
            .in1(N__46604),
            .in2(_gnd_net_),
            .in3(N__46588),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MAIN
