-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 14 2025 21:01:10

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    T01 : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__50557\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50519\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50373\ : std_logic;
signal \N__50370\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50228\ : std_logic;
signal \N__50225\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50139\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50133\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50112\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50103\ : std_logic;
signal \N__50102\ : std_logic;
signal \N__50099\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50062\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50018\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49983\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49976\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49972\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49969\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49966\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49960\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49954\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49938\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49898\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49895\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49892\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49870\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49862\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49859\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49853\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49584\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49559\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49544\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49529\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49511\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49490\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49478\ : std_logic;
signal \N__49475\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49472\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48983\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48963\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48952\ : std_logic;
signal \N__48951\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48929\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48912\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48847\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48540\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48499\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48379\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48246\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48019\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47965\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47952\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47186\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47168\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45985\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45320\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44377\ : std_logic;
signal \N__44374\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44290\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41732\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41681\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41392\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \N_42_i_i\ : std_logic;
signal un7_start_stop_0_a2 : std_logic;
signal \bfn_2_5_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10_cascade_\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_3_7_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_3_8_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal \bfn_3_10_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_149\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31\ : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_154\ : std_logic;
signal pwm_duty_input_2 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_53_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_155\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal il_max_comp2_c : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_153\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_53\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_7_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_72_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_8_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_8_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal il_min_comp1_c : std_logic;
signal il_max_comp1_c : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_enablelt3_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_71\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal s3_phy_c : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal s4_phy_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_397_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_10_25_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_7\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un13_integrator_cry_30\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_26\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.N_166_i_g\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_399_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_i_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.N_1474_i\ : std_logic;
signal \current_shift_inst.control_input_18\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.control_input_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIRB3CP1_0_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.N_54\ : std_logic;
signal \current_shift_inst.timer_s1.N_167_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\ : std_logic;
signal \bfn_13_4_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_8\ : std_logic;
signal \bfn_13_5_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\ : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \elapsed_time_ns_1_RNIPKKEE1_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIOJKEE1_0_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_330_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIRB3CP1_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIJEKEE1_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_286\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_328_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIP93CP1_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNIP93CP1_0_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_310\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal state_ns_i_a2_1 : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \T45_c\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal s1_phy_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \T23_c\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_166_i\ : std_logic;
signal s2_phy_c : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_i_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\ : std_logic;
signal \elapsed_time_ns_1_RNIP7HF91_0_10_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIFJ2591_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIGK2591_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df26\ : std_logic;
signal \elapsed_time_ns_1_RNIOJKEE1_0_7\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal state_3 : std_logic;
signal \T01_c\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_74\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI2IIF91_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI1HIF91_0_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNISBIF91_0_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI0GIF91_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNIP7HF91_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNIQ8HF91_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIR9HF91_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNISAHF91_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNIUCHF91_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_244\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_386_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\ : std_logic;
signal \elapsed_time_ns_1_RNIAE2591_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNII6NQL1_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNII6NQL1_0_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \elapsed_time_ns_1_RNI4HV8E1_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNILGKEE1_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNILGKEE1_0_4_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNI4GU8E1_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNICOU8E1_0_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_397_i_g\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_398_i\ : std_logic;
signal \elapsed_time_ns_1_RNIQ9IF91_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNIRAIF91_0_21\ : std_logic;
signal \elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI3JIF91_0_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23\ : std_logic;
signal \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNIUDIF91_0_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_379_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr9_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIRBJF91_0_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_358\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_354\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIK8NQL1_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6\ : std_logic;
signal \elapsed_time_ns_1_RNINBNQL1_0_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_353\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_353_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_382\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\ : std_logic;
signal \elapsed_time_ns_1_RNIDH2591_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIA965M1_0_18_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNICG2591_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\ : std_logic;
signal \elapsed_time_ns_1_RNI9865M1_0_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lt31_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14\ : std_logic;
signal \elapsed_time_ns_1_RNI6565M1_0_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_395\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_375\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIQENQL1_0_9\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst2.state_RNIG7JFZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI8765M1_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI9865M1_0_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNIBA65M1_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \elapsed_time_ns_1_RNISCJF91_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNIA965M1_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI4FT8E1_0_12_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_369_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_367_clk_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI3FU8E1_0_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \elapsed_time_ns_1_RNIMHKEE1_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_330\ : std_logic;
signal \elapsed_time_ns_1_RNIMHKEE1_0_5_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_328\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \elapsed_time_ns_1_RNIAMU8E1_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNI9LU8E1_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNIBNU8E1_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI8KU8E1_0_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNI5HU8E1_0_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI7JU8E1_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNI6IU8E1_0_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_369\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_344_i_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIGGC6P1_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNIGGC6P1_0_17_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \elapsed_time_ns_1_RNIFFC6P1_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNIIIC6P1_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_318_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \elapsed_time_ns_1_RNIHHC6P1_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \elapsed_time_ns_1_RNI2DT8E1_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \elapsed_time_ns_1_RNI3ET8E1_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \elapsed_time_ns_1_RNI4FT8E1_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_400_i\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst1.N_55\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_RNOZ0Z_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \elapsed_time_ns_1_RNI5GT8E1_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_344_i\ : std_logic;
signal \elapsed_time_ns_1_RNIUE3CP1_0_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \elapsed_time_ns_1_RNI7IT8E1_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_269_iZ0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNI7IT8E1_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \elapsed_time_ns_1_RNI1I3CP1_0_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_367_clk\ : std_logic;
signal \delay_measurement_inst.delay_tr9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \elapsed_time_ns_1_RNI5IV8E1_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.N_318\ : std_logic;
signal \elapsed_time_ns_1_RNIDDC6P1_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \T12_c\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_399_i_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_394\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_346\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_346_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_349\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_349_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_351\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_362\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_362_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\ : std_logic;
signal \delay_measurement_inst.N_365\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21354\&\N__21347\&\N__21352\&\N__21346\&\N__21353\&\N__21345\&\N__21355\&\N__21342\&\N__21348\&\N__21341\&\N__21349\&\N__21343\&\N__21350\&\N__21344\&\N__21351\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28313\&\N__28303\&'0'&'0'&'0'&\N__28301\&\N__28312\&\N__28302\&\N__28311\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__21406\&\N__21409\&\N__21407\&\N__21410\&\N__21408\&\N__21914\&\N__21839\&\N__21722\&\N__21878\&\N__21690\&\N__21644\&\N__22390\&\N__21745\&\N__20257\&\N__20242\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28288\&\N__28285\&'0'&'0'&'0'&\N__28283\&\N__28287\&\N__28284\&\N__28286\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__21169\,
            RESETB => \N__34198\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__28314\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__28300\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__28289\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__28282\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__50555\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50557\,
            DIN => \N__50556\,
            DOUT => \N__50555\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50557\,
            PADOUT => \N__50556\,
            PADIN => \N__50555\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50546\,
            DIN => \N__50545\,
            DOUT => \N__50544\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50546\,
            PADOUT => \N__50545\,
            PADIN => \N__50544\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__38215\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50537\,
            DIN => \N__50536\,
            DOUT => \N__50535\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50537\,
            PADOUT => \N__50536\,
            PADIN => \N__50535\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50528\,
            DIN => \N__50527\,
            DOUT => \N__50526\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50528\,
            PADOUT => \N__50527\,
            PADIN => \N__50526\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50519\,
            DIN => \N__50518\,
            DOUT => \N__50517\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50519\,
            PADOUT => \N__50518\,
            PADIN => \N__50517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34900\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50510\,
            DIN => \N__50509\,
            DOUT => \N__50508\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50510\,
            PADOUT => \N__50509\,
            PADIN => \N__50508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20896\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50501\,
            DIN => \N__50500\,
            DOUT => \N__50499\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50501\,
            PADOUT => \N__50500\,
            PADIN => \N__50499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50492\,
            DIN => \N__50491\,
            DOUT => \N__50490\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50492\,
            PADOUT => \N__50491\,
            PADIN => \N__50490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34822\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50483\,
            DIN => \N__50482\,
            DOUT => \N__50481\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50483\,
            PADOUT => \N__50482\,
            PADIN => \N__50481\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__46555\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50474\,
            DIN => \N__50473\,
            DOUT => \N__50472\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50474\,
            PADOUT => \N__50473\,
            PADIN => \N__50472\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50465\,
            DIN => \N__50464\,
            DOUT => \N__50463\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50465\,
            PADOUT => \N__50464\,
            PADIN => \N__50463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34942\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50456\,
            DIN => \N__50455\,
            DOUT => \N__50454\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50456\,
            PADOUT => \N__50455\,
            PADIN => \N__50454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50447\,
            DIN => \N__50446\,
            DOUT => \N__50445\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50447\,
            PADOUT => \N__50446\,
            PADIN => \N__50445\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50438\,
            DIN => \N__50437\,
            DOUT => \N__50436\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50438\,
            PADOUT => \N__50437\,
            PADIN => \N__50436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25132\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50429\,
            DIN => \N__50428\,
            DOUT => \N__50427\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50429\,
            PADOUT => \N__50428\,
            PADIN => \N__50427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34630\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50420\,
            DIN => \N__50419\,
            DOUT => \N__50418\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50420\,
            PADOUT => \N__50419\,
            PADIN => \N__50418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50411\,
            DIN => \N__50410\,
            DOUT => \N__50409\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50411\,
            PADOUT => \N__50410\,
            PADIN => \N__50409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11955\ : InMux
    port map (
            O => \N__50392\,
            I => \N__50388\
        );

    \I__11954\ : InMux
    port map (
            O => \N__50391\,
            I => \N__50385\
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__50388\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__50385\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__11951\ : InMux
    port map (
            O => \N__50380\,
            I => \N__50376\
        );

    \I__11950\ : InMux
    port map (
            O => \N__50379\,
            I => \N__50373\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__50376\,
            I => \N__50370\
        );

    \I__11948\ : LocalMux
    port map (
            O => \N__50373\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__11947\ : Odrv4
    port map (
            O => \N__50370\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__11946\ : InMux
    port map (
            O => \N__50365\,
            I => \N__50362\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__50362\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df24\
        );

    \I__11944\ : InMux
    port map (
            O => \N__50359\,
            I => \N__50355\
        );

    \I__11943\ : InMux
    port map (
            O => \N__50358\,
            I => \N__50352\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__50355\,
            I => \N__50349\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__50352\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__11940\ : Odrv4
    port map (
            O => \N__50349\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__11939\ : InMux
    port map (
            O => \N__50344\,
            I => \N__50340\
        );

    \I__11938\ : InMux
    port map (
            O => \N__50343\,
            I => \N__50337\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__50340\,
            I => \N__50334\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__50337\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__11935\ : Odrv4
    port map (
            O => \N__50334\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__11934\ : InMux
    port map (
            O => \N__50329\,
            I => \N__50326\
        );

    \I__11933\ : LocalMux
    port map (
            O => \N__50326\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df20\
        );

    \I__11932\ : CEMux
    port map (
            O => \N__50323\,
            I => \N__50317\
        );

    \I__11931\ : CEMux
    port map (
            O => \N__50322\,
            I => \N__50314\
        );

    \I__11930\ : CEMux
    port map (
            O => \N__50321\,
            I => \N__50311\
        );

    \I__11929\ : CEMux
    port map (
            O => \N__50320\,
            I => \N__50308\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__50317\,
            I => \N__50296\
        );

    \I__11927\ : LocalMux
    port map (
            O => \N__50314\,
            I => \N__50296\
        );

    \I__11926\ : LocalMux
    port map (
            O => \N__50311\,
            I => \N__50285\
        );

    \I__11925\ : LocalMux
    port map (
            O => \N__50308\,
            I => \N__50266\
        );

    \I__11924\ : InMux
    port map (
            O => \N__50307\,
            I => \N__50259\
        );

    \I__11923\ : InMux
    port map (
            O => \N__50306\,
            I => \N__50259\
        );

    \I__11922\ : InMux
    port map (
            O => \N__50305\,
            I => \N__50259\
        );

    \I__11921\ : InMux
    port map (
            O => \N__50304\,
            I => \N__50250\
        );

    \I__11920\ : InMux
    port map (
            O => \N__50303\,
            I => \N__50250\
        );

    \I__11919\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50250\
        );

    \I__11918\ : InMux
    port map (
            O => \N__50301\,
            I => \N__50250\
        );

    \I__11917\ : Span4Mux_v
    port map (
            O => \N__50296\,
            I => \N__50247\
        );

    \I__11916\ : InMux
    port map (
            O => \N__50295\,
            I => \N__50240\
        );

    \I__11915\ : InMux
    port map (
            O => \N__50294\,
            I => \N__50240\
        );

    \I__11914\ : InMux
    port map (
            O => \N__50293\,
            I => \N__50240\
        );

    \I__11913\ : InMux
    port map (
            O => \N__50292\,
            I => \N__50237\
        );

    \I__11912\ : InMux
    port map (
            O => \N__50291\,
            I => \N__50228\
        );

    \I__11911\ : InMux
    port map (
            O => \N__50290\,
            I => \N__50228\
        );

    \I__11910\ : InMux
    port map (
            O => \N__50289\,
            I => \N__50228\
        );

    \I__11909\ : InMux
    port map (
            O => \N__50288\,
            I => \N__50228\
        );

    \I__11908\ : Span4Mux_v
    port map (
            O => \N__50285\,
            I => \N__50225\
        );

    \I__11907\ : InMux
    port map (
            O => \N__50284\,
            I => \N__50216\
        );

    \I__11906\ : InMux
    port map (
            O => \N__50283\,
            I => \N__50216\
        );

    \I__11905\ : InMux
    port map (
            O => \N__50282\,
            I => \N__50216\
        );

    \I__11904\ : InMux
    port map (
            O => \N__50281\,
            I => \N__50216\
        );

    \I__11903\ : InMux
    port map (
            O => \N__50280\,
            I => \N__50207\
        );

    \I__11902\ : InMux
    port map (
            O => \N__50279\,
            I => \N__50207\
        );

    \I__11901\ : InMux
    port map (
            O => \N__50278\,
            I => \N__50207\
        );

    \I__11900\ : InMux
    port map (
            O => \N__50277\,
            I => \N__50207\
        );

    \I__11899\ : InMux
    port map (
            O => \N__50276\,
            I => \N__50198\
        );

    \I__11898\ : InMux
    port map (
            O => \N__50275\,
            I => \N__50198\
        );

    \I__11897\ : InMux
    port map (
            O => \N__50274\,
            I => \N__50198\
        );

    \I__11896\ : InMux
    port map (
            O => \N__50273\,
            I => \N__50198\
        );

    \I__11895\ : InMux
    port map (
            O => \N__50272\,
            I => \N__50189\
        );

    \I__11894\ : InMux
    port map (
            O => \N__50271\,
            I => \N__50189\
        );

    \I__11893\ : InMux
    port map (
            O => \N__50270\,
            I => \N__50189\
        );

    \I__11892\ : InMux
    port map (
            O => \N__50269\,
            I => \N__50189\
        );

    \I__11891\ : Span4Mux_v
    port map (
            O => \N__50266\,
            I => \N__50184\
        );

    \I__11890\ : LocalMux
    port map (
            O => \N__50259\,
            I => \N__50184\
        );

    \I__11889\ : LocalMux
    port map (
            O => \N__50250\,
            I => \N__50181\
        );

    \I__11888\ : Span4Mux_h
    port map (
            O => \N__50247\,
            I => \N__50172\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__50240\,
            I => \N__50172\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__50237\,
            I => \N__50172\
        );

    \I__11885\ : LocalMux
    port map (
            O => \N__50228\,
            I => \N__50172\
        );

    \I__11884\ : Span4Mux_h
    port map (
            O => \N__50225\,
            I => \N__50165\
        );

    \I__11883\ : LocalMux
    port map (
            O => \N__50216\,
            I => \N__50165\
        );

    \I__11882\ : LocalMux
    port map (
            O => \N__50207\,
            I => \N__50165\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__50198\,
            I => \N__50160\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__50189\,
            I => \N__50160\
        );

    \I__11879\ : Span4Mux_h
    port map (
            O => \N__50184\,
            I => \N__50155\
        );

    \I__11878\ : Span4Mux_h
    port map (
            O => \N__50181\,
            I => \N__50155\
        );

    \I__11877\ : Span4Mux_h
    port map (
            O => \N__50172\,
            I => \N__50152\
        );

    \I__11876\ : Span4Mux_h
    port map (
            O => \N__50165\,
            I => \N__50149\
        );

    \I__11875\ : Odrv4
    port map (
            O => \N__50160\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11874\ : Odrv4
    port map (
            O => \N__50155\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11873\ : Odrv4
    port map (
            O => \N__50152\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11872\ : Odrv4
    port map (
            O => \N__50149\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11871\ : InMux
    port map (
            O => \N__50140\,
            I => \N__50136\
        );

    \I__11870\ : InMux
    port map (
            O => \N__50139\,
            I => \N__50133\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__50136\,
            I => \N__50128\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__50133\,
            I => \N__50125\
        );

    \I__11867\ : InMux
    port map (
            O => \N__50132\,
            I => \N__50122\
        );

    \I__11866\ : InMux
    port map (
            O => \N__50131\,
            I => \N__50119\
        );

    \I__11865\ : Span4Mux_v
    port map (
            O => \N__50128\,
            I => \N__50112\
        );

    \I__11864\ : Span4Mux_v
    port map (
            O => \N__50125\,
            I => \N__50112\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__50122\,
            I => \N__50112\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__50119\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11861\ : Odrv4
    port map (
            O => \N__50112\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11860\ : InMux
    port map (
            O => \N__50107\,
            I => \N__50103\
        );

    \I__11859\ : InMux
    port map (
            O => \N__50106\,
            I => \N__50099\
        );

    \I__11858\ : LocalMux
    port map (
            O => \N__50103\,
            I => \N__50095\
        );

    \I__11857\ : InMux
    port map (
            O => \N__50102\,
            I => \N__50092\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__50099\,
            I => \N__50089\
        );

    \I__11855\ : InMux
    port map (
            O => \N__50098\,
            I => \N__50085\
        );

    \I__11854\ : Span12Mux_h
    port map (
            O => \N__50095\,
            I => \N__50082\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__50092\,
            I => \N__50079\
        );

    \I__11852\ : Span4Mux_v
    port map (
            O => \N__50089\,
            I => \N__50076\
        );

    \I__11851\ : InMux
    port map (
            O => \N__50088\,
            I => \N__50073\
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__50085\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__11849\ : Odrv12
    port map (
            O => \N__50082\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__11848\ : Odrv4
    port map (
            O => \N__50079\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__11847\ : Odrv4
    port map (
            O => \N__50076\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__50073\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__11845\ : InMux
    port map (
            O => \N__50062\,
            I => \N__50059\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__50059\,
            I => \N__50055\
        );

    \I__11843\ : InMux
    port map (
            O => \N__50058\,
            I => \N__50052\
        );

    \I__11842\ : Span4Mux_h
    port map (
            O => \N__50055\,
            I => \N__50049\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__50052\,
            I => \N__50046\
        );

    \I__11840\ : Span4Mux_h
    port map (
            O => \N__50049\,
            I => \N__50041\
        );

    \I__11839\ : Span4Mux_h
    port map (
            O => \N__50046\,
            I => \N__50041\
        );

    \I__11838\ : Odrv4
    port map (
            O => \N__50041\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__11837\ : CascadeMux
    port map (
            O => \N__50038\,
            I => \N__50034\
        );

    \I__11836\ : CascadeMux
    port map (
            O => \N__50037\,
            I => \N__50031\
        );

    \I__11835\ : InMux
    port map (
            O => \N__50034\,
            I => \N__50028\
        );

    \I__11834\ : InMux
    port map (
            O => \N__50031\,
            I => \N__50025\
        );

    \I__11833\ : LocalMux
    port map (
            O => \N__50028\,
            I => \N__50022\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__50025\,
            I => \N__50019\
        );

    \I__11831\ : Span4Mux_v
    port map (
            O => \N__50022\,
            I => \N__50011\
        );

    \I__11830\ : Span4Mux_v
    port map (
            O => \N__50019\,
            I => \N__50011\
        );

    \I__11829\ : InMux
    port map (
            O => \N__50018\,
            I => \N__50006\
        );

    \I__11828\ : InMux
    port map (
            O => \N__50017\,
            I => \N__50006\
        );

    \I__11827\ : InMux
    port map (
            O => \N__50016\,
            I => \N__50003\
        );

    \I__11826\ : Sp12to4
    port map (
            O => \N__50011\,
            I => \N__49998\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__50006\,
            I => \N__49998\
        );

    \I__11824\ : LocalMux
    port map (
            O => \N__50003\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__11823\ : Odrv12
    port map (
            O => \N__49998\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__11822\ : CascadeMux
    port map (
            O => \N__49993\,
            I => \N__49990\
        );

    \I__11821\ : InMux
    port map (
            O => \N__49990\,
            I => \N__49986\
        );

    \I__11820\ : InMux
    port map (
            O => \N__49989\,
            I => \N__49983\
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__49986\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__11818\ : LocalMux
    port map (
            O => \N__49983\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__11817\ : ClkMux
    port map (
            O => \N__49978\,
            I => \N__49591\
        );

    \I__11816\ : ClkMux
    port map (
            O => \N__49977\,
            I => \N__49591\
        );

    \I__11815\ : ClkMux
    port map (
            O => \N__49976\,
            I => \N__49591\
        );

    \I__11814\ : ClkMux
    port map (
            O => \N__49975\,
            I => \N__49591\
        );

    \I__11813\ : ClkMux
    port map (
            O => \N__49974\,
            I => \N__49591\
        );

    \I__11812\ : ClkMux
    port map (
            O => \N__49973\,
            I => \N__49591\
        );

    \I__11811\ : ClkMux
    port map (
            O => \N__49972\,
            I => \N__49591\
        );

    \I__11810\ : ClkMux
    port map (
            O => \N__49971\,
            I => \N__49591\
        );

    \I__11809\ : ClkMux
    port map (
            O => \N__49970\,
            I => \N__49591\
        );

    \I__11808\ : ClkMux
    port map (
            O => \N__49969\,
            I => \N__49591\
        );

    \I__11807\ : ClkMux
    port map (
            O => \N__49968\,
            I => \N__49591\
        );

    \I__11806\ : ClkMux
    port map (
            O => \N__49967\,
            I => \N__49591\
        );

    \I__11805\ : ClkMux
    port map (
            O => \N__49966\,
            I => \N__49591\
        );

    \I__11804\ : ClkMux
    port map (
            O => \N__49965\,
            I => \N__49591\
        );

    \I__11803\ : ClkMux
    port map (
            O => \N__49964\,
            I => \N__49591\
        );

    \I__11802\ : ClkMux
    port map (
            O => \N__49963\,
            I => \N__49591\
        );

    \I__11801\ : ClkMux
    port map (
            O => \N__49962\,
            I => \N__49591\
        );

    \I__11800\ : ClkMux
    port map (
            O => \N__49961\,
            I => \N__49591\
        );

    \I__11799\ : ClkMux
    port map (
            O => \N__49960\,
            I => \N__49591\
        );

    \I__11798\ : ClkMux
    port map (
            O => \N__49959\,
            I => \N__49591\
        );

    \I__11797\ : ClkMux
    port map (
            O => \N__49958\,
            I => \N__49591\
        );

    \I__11796\ : ClkMux
    port map (
            O => \N__49957\,
            I => \N__49591\
        );

    \I__11795\ : ClkMux
    port map (
            O => \N__49956\,
            I => \N__49591\
        );

    \I__11794\ : ClkMux
    port map (
            O => \N__49955\,
            I => \N__49591\
        );

    \I__11793\ : ClkMux
    port map (
            O => \N__49954\,
            I => \N__49591\
        );

    \I__11792\ : ClkMux
    port map (
            O => \N__49953\,
            I => \N__49591\
        );

    \I__11791\ : ClkMux
    port map (
            O => \N__49952\,
            I => \N__49591\
        );

    \I__11790\ : ClkMux
    port map (
            O => \N__49951\,
            I => \N__49591\
        );

    \I__11789\ : ClkMux
    port map (
            O => \N__49950\,
            I => \N__49591\
        );

    \I__11788\ : ClkMux
    port map (
            O => \N__49949\,
            I => \N__49591\
        );

    \I__11787\ : ClkMux
    port map (
            O => \N__49948\,
            I => \N__49591\
        );

    \I__11786\ : ClkMux
    port map (
            O => \N__49947\,
            I => \N__49591\
        );

    \I__11785\ : ClkMux
    port map (
            O => \N__49946\,
            I => \N__49591\
        );

    \I__11784\ : ClkMux
    port map (
            O => \N__49945\,
            I => \N__49591\
        );

    \I__11783\ : ClkMux
    port map (
            O => \N__49944\,
            I => \N__49591\
        );

    \I__11782\ : ClkMux
    port map (
            O => \N__49943\,
            I => \N__49591\
        );

    \I__11781\ : ClkMux
    port map (
            O => \N__49942\,
            I => \N__49591\
        );

    \I__11780\ : ClkMux
    port map (
            O => \N__49941\,
            I => \N__49591\
        );

    \I__11779\ : ClkMux
    port map (
            O => \N__49940\,
            I => \N__49591\
        );

    \I__11778\ : ClkMux
    port map (
            O => \N__49939\,
            I => \N__49591\
        );

    \I__11777\ : ClkMux
    port map (
            O => \N__49938\,
            I => \N__49591\
        );

    \I__11776\ : ClkMux
    port map (
            O => \N__49937\,
            I => \N__49591\
        );

    \I__11775\ : ClkMux
    port map (
            O => \N__49936\,
            I => \N__49591\
        );

    \I__11774\ : ClkMux
    port map (
            O => \N__49935\,
            I => \N__49591\
        );

    \I__11773\ : ClkMux
    port map (
            O => \N__49934\,
            I => \N__49591\
        );

    \I__11772\ : ClkMux
    port map (
            O => \N__49933\,
            I => \N__49591\
        );

    \I__11771\ : ClkMux
    port map (
            O => \N__49932\,
            I => \N__49591\
        );

    \I__11770\ : ClkMux
    port map (
            O => \N__49931\,
            I => \N__49591\
        );

    \I__11769\ : ClkMux
    port map (
            O => \N__49930\,
            I => \N__49591\
        );

    \I__11768\ : ClkMux
    port map (
            O => \N__49929\,
            I => \N__49591\
        );

    \I__11767\ : ClkMux
    port map (
            O => \N__49928\,
            I => \N__49591\
        );

    \I__11766\ : ClkMux
    port map (
            O => \N__49927\,
            I => \N__49591\
        );

    \I__11765\ : ClkMux
    port map (
            O => \N__49926\,
            I => \N__49591\
        );

    \I__11764\ : ClkMux
    port map (
            O => \N__49925\,
            I => \N__49591\
        );

    \I__11763\ : ClkMux
    port map (
            O => \N__49924\,
            I => \N__49591\
        );

    \I__11762\ : ClkMux
    port map (
            O => \N__49923\,
            I => \N__49591\
        );

    \I__11761\ : ClkMux
    port map (
            O => \N__49922\,
            I => \N__49591\
        );

    \I__11760\ : ClkMux
    port map (
            O => \N__49921\,
            I => \N__49591\
        );

    \I__11759\ : ClkMux
    port map (
            O => \N__49920\,
            I => \N__49591\
        );

    \I__11758\ : ClkMux
    port map (
            O => \N__49919\,
            I => \N__49591\
        );

    \I__11757\ : ClkMux
    port map (
            O => \N__49918\,
            I => \N__49591\
        );

    \I__11756\ : ClkMux
    port map (
            O => \N__49917\,
            I => \N__49591\
        );

    \I__11755\ : ClkMux
    port map (
            O => \N__49916\,
            I => \N__49591\
        );

    \I__11754\ : ClkMux
    port map (
            O => \N__49915\,
            I => \N__49591\
        );

    \I__11753\ : ClkMux
    port map (
            O => \N__49914\,
            I => \N__49591\
        );

    \I__11752\ : ClkMux
    port map (
            O => \N__49913\,
            I => \N__49591\
        );

    \I__11751\ : ClkMux
    port map (
            O => \N__49912\,
            I => \N__49591\
        );

    \I__11750\ : ClkMux
    port map (
            O => \N__49911\,
            I => \N__49591\
        );

    \I__11749\ : ClkMux
    port map (
            O => \N__49910\,
            I => \N__49591\
        );

    \I__11748\ : ClkMux
    port map (
            O => \N__49909\,
            I => \N__49591\
        );

    \I__11747\ : ClkMux
    port map (
            O => \N__49908\,
            I => \N__49591\
        );

    \I__11746\ : ClkMux
    port map (
            O => \N__49907\,
            I => \N__49591\
        );

    \I__11745\ : ClkMux
    port map (
            O => \N__49906\,
            I => \N__49591\
        );

    \I__11744\ : ClkMux
    port map (
            O => \N__49905\,
            I => \N__49591\
        );

    \I__11743\ : ClkMux
    port map (
            O => \N__49904\,
            I => \N__49591\
        );

    \I__11742\ : ClkMux
    port map (
            O => \N__49903\,
            I => \N__49591\
        );

    \I__11741\ : ClkMux
    port map (
            O => \N__49902\,
            I => \N__49591\
        );

    \I__11740\ : ClkMux
    port map (
            O => \N__49901\,
            I => \N__49591\
        );

    \I__11739\ : ClkMux
    port map (
            O => \N__49900\,
            I => \N__49591\
        );

    \I__11738\ : ClkMux
    port map (
            O => \N__49899\,
            I => \N__49591\
        );

    \I__11737\ : ClkMux
    port map (
            O => \N__49898\,
            I => \N__49591\
        );

    \I__11736\ : ClkMux
    port map (
            O => \N__49897\,
            I => \N__49591\
        );

    \I__11735\ : ClkMux
    port map (
            O => \N__49896\,
            I => \N__49591\
        );

    \I__11734\ : ClkMux
    port map (
            O => \N__49895\,
            I => \N__49591\
        );

    \I__11733\ : ClkMux
    port map (
            O => \N__49894\,
            I => \N__49591\
        );

    \I__11732\ : ClkMux
    port map (
            O => \N__49893\,
            I => \N__49591\
        );

    \I__11731\ : ClkMux
    port map (
            O => \N__49892\,
            I => \N__49591\
        );

    \I__11730\ : ClkMux
    port map (
            O => \N__49891\,
            I => \N__49591\
        );

    \I__11729\ : ClkMux
    port map (
            O => \N__49890\,
            I => \N__49591\
        );

    \I__11728\ : ClkMux
    port map (
            O => \N__49889\,
            I => \N__49591\
        );

    \I__11727\ : ClkMux
    port map (
            O => \N__49888\,
            I => \N__49591\
        );

    \I__11726\ : ClkMux
    port map (
            O => \N__49887\,
            I => \N__49591\
        );

    \I__11725\ : ClkMux
    port map (
            O => \N__49886\,
            I => \N__49591\
        );

    \I__11724\ : ClkMux
    port map (
            O => \N__49885\,
            I => \N__49591\
        );

    \I__11723\ : ClkMux
    port map (
            O => \N__49884\,
            I => \N__49591\
        );

    \I__11722\ : ClkMux
    port map (
            O => \N__49883\,
            I => \N__49591\
        );

    \I__11721\ : ClkMux
    port map (
            O => \N__49882\,
            I => \N__49591\
        );

    \I__11720\ : ClkMux
    port map (
            O => \N__49881\,
            I => \N__49591\
        );

    \I__11719\ : ClkMux
    port map (
            O => \N__49880\,
            I => \N__49591\
        );

    \I__11718\ : ClkMux
    port map (
            O => \N__49879\,
            I => \N__49591\
        );

    \I__11717\ : ClkMux
    port map (
            O => \N__49878\,
            I => \N__49591\
        );

    \I__11716\ : ClkMux
    port map (
            O => \N__49877\,
            I => \N__49591\
        );

    \I__11715\ : ClkMux
    port map (
            O => \N__49876\,
            I => \N__49591\
        );

    \I__11714\ : ClkMux
    port map (
            O => \N__49875\,
            I => \N__49591\
        );

    \I__11713\ : ClkMux
    port map (
            O => \N__49874\,
            I => \N__49591\
        );

    \I__11712\ : ClkMux
    port map (
            O => \N__49873\,
            I => \N__49591\
        );

    \I__11711\ : ClkMux
    port map (
            O => \N__49872\,
            I => \N__49591\
        );

    \I__11710\ : ClkMux
    port map (
            O => \N__49871\,
            I => \N__49591\
        );

    \I__11709\ : ClkMux
    port map (
            O => \N__49870\,
            I => \N__49591\
        );

    \I__11708\ : ClkMux
    port map (
            O => \N__49869\,
            I => \N__49591\
        );

    \I__11707\ : ClkMux
    port map (
            O => \N__49868\,
            I => \N__49591\
        );

    \I__11706\ : ClkMux
    port map (
            O => \N__49867\,
            I => \N__49591\
        );

    \I__11705\ : ClkMux
    port map (
            O => \N__49866\,
            I => \N__49591\
        );

    \I__11704\ : ClkMux
    port map (
            O => \N__49865\,
            I => \N__49591\
        );

    \I__11703\ : ClkMux
    port map (
            O => \N__49864\,
            I => \N__49591\
        );

    \I__11702\ : ClkMux
    port map (
            O => \N__49863\,
            I => \N__49591\
        );

    \I__11701\ : ClkMux
    port map (
            O => \N__49862\,
            I => \N__49591\
        );

    \I__11700\ : ClkMux
    port map (
            O => \N__49861\,
            I => \N__49591\
        );

    \I__11699\ : ClkMux
    port map (
            O => \N__49860\,
            I => \N__49591\
        );

    \I__11698\ : ClkMux
    port map (
            O => \N__49859\,
            I => \N__49591\
        );

    \I__11697\ : ClkMux
    port map (
            O => \N__49858\,
            I => \N__49591\
        );

    \I__11696\ : ClkMux
    port map (
            O => \N__49857\,
            I => \N__49591\
        );

    \I__11695\ : ClkMux
    port map (
            O => \N__49856\,
            I => \N__49591\
        );

    \I__11694\ : ClkMux
    port map (
            O => \N__49855\,
            I => \N__49591\
        );

    \I__11693\ : ClkMux
    port map (
            O => \N__49854\,
            I => \N__49591\
        );

    \I__11692\ : ClkMux
    port map (
            O => \N__49853\,
            I => \N__49591\
        );

    \I__11691\ : ClkMux
    port map (
            O => \N__49852\,
            I => \N__49591\
        );

    \I__11690\ : ClkMux
    port map (
            O => \N__49851\,
            I => \N__49591\
        );

    \I__11689\ : ClkMux
    port map (
            O => \N__49850\,
            I => \N__49591\
        );

    \I__11688\ : GlobalMux
    port map (
            O => \N__49591\,
            I => clk_100mhz_0
        );

    \I__11687\ : InMux
    port map (
            O => \N__49588\,
            I => \N__49577\
        );

    \I__11686\ : InMux
    port map (
            O => \N__49587\,
            I => \N__49574\
        );

    \I__11685\ : InMux
    port map (
            O => \N__49586\,
            I => \N__49571\
        );

    \I__11684\ : InMux
    port map (
            O => \N__49585\,
            I => \N__49568\
        );

    \I__11683\ : InMux
    port map (
            O => \N__49584\,
            I => \N__49565\
        );

    \I__11682\ : InMux
    port map (
            O => \N__49583\,
            I => \N__49562\
        );

    \I__11681\ : InMux
    port map (
            O => \N__49582\,
            I => \N__49559\
        );

    \I__11680\ : InMux
    port map (
            O => \N__49581\,
            I => \N__49554\
        );

    \I__11679\ : InMux
    port map (
            O => \N__49580\,
            I => \N__49554\
        );

    \I__11678\ : LocalMux
    port map (
            O => \N__49577\,
            I => \N__49551\
        );

    \I__11677\ : LocalMux
    port map (
            O => \N__49574\,
            I => \N__49548\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__49571\,
            I => \N__49545\
        );

    \I__11675\ : LocalMux
    port map (
            O => \N__49568\,
            I => \N__49475\
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__49565\,
            I => \N__49453\
        );

    \I__11673\ : LocalMux
    port map (
            O => \N__49562\,
            I => \N__49445\
        );

    \I__11672\ : LocalMux
    port map (
            O => \N__49559\,
            I => \N__49427\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__49554\,
            I => \N__49417\
        );

    \I__11670\ : Glb2LocalMux
    port map (
            O => \N__49551\,
            I => \N__49138\
        );

    \I__11669\ : Glb2LocalMux
    port map (
            O => \N__49548\,
            I => \N__49138\
        );

    \I__11668\ : Glb2LocalMux
    port map (
            O => \N__49545\,
            I => \N__49138\
        );

    \I__11667\ : SRMux
    port map (
            O => \N__49544\,
            I => \N__49138\
        );

    \I__11666\ : SRMux
    port map (
            O => \N__49543\,
            I => \N__49138\
        );

    \I__11665\ : SRMux
    port map (
            O => \N__49542\,
            I => \N__49138\
        );

    \I__11664\ : SRMux
    port map (
            O => \N__49541\,
            I => \N__49138\
        );

    \I__11663\ : SRMux
    port map (
            O => \N__49540\,
            I => \N__49138\
        );

    \I__11662\ : SRMux
    port map (
            O => \N__49539\,
            I => \N__49138\
        );

    \I__11661\ : SRMux
    port map (
            O => \N__49538\,
            I => \N__49138\
        );

    \I__11660\ : SRMux
    port map (
            O => \N__49537\,
            I => \N__49138\
        );

    \I__11659\ : SRMux
    port map (
            O => \N__49536\,
            I => \N__49138\
        );

    \I__11658\ : SRMux
    port map (
            O => \N__49535\,
            I => \N__49138\
        );

    \I__11657\ : SRMux
    port map (
            O => \N__49534\,
            I => \N__49138\
        );

    \I__11656\ : SRMux
    port map (
            O => \N__49533\,
            I => \N__49138\
        );

    \I__11655\ : SRMux
    port map (
            O => \N__49532\,
            I => \N__49138\
        );

    \I__11654\ : SRMux
    port map (
            O => \N__49531\,
            I => \N__49138\
        );

    \I__11653\ : SRMux
    port map (
            O => \N__49530\,
            I => \N__49138\
        );

    \I__11652\ : SRMux
    port map (
            O => \N__49529\,
            I => \N__49138\
        );

    \I__11651\ : SRMux
    port map (
            O => \N__49528\,
            I => \N__49138\
        );

    \I__11650\ : SRMux
    port map (
            O => \N__49527\,
            I => \N__49138\
        );

    \I__11649\ : SRMux
    port map (
            O => \N__49526\,
            I => \N__49138\
        );

    \I__11648\ : SRMux
    port map (
            O => \N__49525\,
            I => \N__49138\
        );

    \I__11647\ : SRMux
    port map (
            O => \N__49524\,
            I => \N__49138\
        );

    \I__11646\ : SRMux
    port map (
            O => \N__49523\,
            I => \N__49138\
        );

    \I__11645\ : SRMux
    port map (
            O => \N__49522\,
            I => \N__49138\
        );

    \I__11644\ : SRMux
    port map (
            O => \N__49521\,
            I => \N__49138\
        );

    \I__11643\ : SRMux
    port map (
            O => \N__49520\,
            I => \N__49138\
        );

    \I__11642\ : SRMux
    port map (
            O => \N__49519\,
            I => \N__49138\
        );

    \I__11641\ : SRMux
    port map (
            O => \N__49518\,
            I => \N__49138\
        );

    \I__11640\ : SRMux
    port map (
            O => \N__49517\,
            I => \N__49138\
        );

    \I__11639\ : SRMux
    port map (
            O => \N__49516\,
            I => \N__49138\
        );

    \I__11638\ : SRMux
    port map (
            O => \N__49515\,
            I => \N__49138\
        );

    \I__11637\ : SRMux
    port map (
            O => \N__49514\,
            I => \N__49138\
        );

    \I__11636\ : SRMux
    port map (
            O => \N__49513\,
            I => \N__49138\
        );

    \I__11635\ : SRMux
    port map (
            O => \N__49512\,
            I => \N__49138\
        );

    \I__11634\ : SRMux
    port map (
            O => \N__49511\,
            I => \N__49138\
        );

    \I__11633\ : SRMux
    port map (
            O => \N__49510\,
            I => \N__49138\
        );

    \I__11632\ : SRMux
    port map (
            O => \N__49509\,
            I => \N__49138\
        );

    \I__11631\ : SRMux
    port map (
            O => \N__49508\,
            I => \N__49138\
        );

    \I__11630\ : SRMux
    port map (
            O => \N__49507\,
            I => \N__49138\
        );

    \I__11629\ : SRMux
    port map (
            O => \N__49506\,
            I => \N__49138\
        );

    \I__11628\ : SRMux
    port map (
            O => \N__49505\,
            I => \N__49138\
        );

    \I__11627\ : SRMux
    port map (
            O => \N__49504\,
            I => \N__49138\
        );

    \I__11626\ : SRMux
    port map (
            O => \N__49503\,
            I => \N__49138\
        );

    \I__11625\ : SRMux
    port map (
            O => \N__49502\,
            I => \N__49138\
        );

    \I__11624\ : SRMux
    port map (
            O => \N__49501\,
            I => \N__49138\
        );

    \I__11623\ : SRMux
    port map (
            O => \N__49500\,
            I => \N__49138\
        );

    \I__11622\ : SRMux
    port map (
            O => \N__49499\,
            I => \N__49138\
        );

    \I__11621\ : SRMux
    port map (
            O => \N__49498\,
            I => \N__49138\
        );

    \I__11620\ : SRMux
    port map (
            O => \N__49497\,
            I => \N__49138\
        );

    \I__11619\ : SRMux
    port map (
            O => \N__49496\,
            I => \N__49138\
        );

    \I__11618\ : SRMux
    port map (
            O => \N__49495\,
            I => \N__49138\
        );

    \I__11617\ : SRMux
    port map (
            O => \N__49494\,
            I => \N__49138\
        );

    \I__11616\ : SRMux
    port map (
            O => \N__49493\,
            I => \N__49138\
        );

    \I__11615\ : SRMux
    port map (
            O => \N__49492\,
            I => \N__49138\
        );

    \I__11614\ : SRMux
    port map (
            O => \N__49491\,
            I => \N__49138\
        );

    \I__11613\ : SRMux
    port map (
            O => \N__49490\,
            I => \N__49138\
        );

    \I__11612\ : SRMux
    port map (
            O => \N__49489\,
            I => \N__49138\
        );

    \I__11611\ : SRMux
    port map (
            O => \N__49488\,
            I => \N__49138\
        );

    \I__11610\ : SRMux
    port map (
            O => \N__49487\,
            I => \N__49138\
        );

    \I__11609\ : SRMux
    port map (
            O => \N__49486\,
            I => \N__49138\
        );

    \I__11608\ : SRMux
    port map (
            O => \N__49485\,
            I => \N__49138\
        );

    \I__11607\ : SRMux
    port map (
            O => \N__49484\,
            I => \N__49138\
        );

    \I__11606\ : SRMux
    port map (
            O => \N__49483\,
            I => \N__49138\
        );

    \I__11605\ : SRMux
    port map (
            O => \N__49482\,
            I => \N__49138\
        );

    \I__11604\ : SRMux
    port map (
            O => \N__49481\,
            I => \N__49138\
        );

    \I__11603\ : SRMux
    port map (
            O => \N__49480\,
            I => \N__49138\
        );

    \I__11602\ : SRMux
    port map (
            O => \N__49479\,
            I => \N__49138\
        );

    \I__11601\ : SRMux
    port map (
            O => \N__49478\,
            I => \N__49138\
        );

    \I__11600\ : Glb2LocalMux
    port map (
            O => \N__49475\,
            I => \N__49138\
        );

    \I__11599\ : SRMux
    port map (
            O => \N__49474\,
            I => \N__49138\
        );

    \I__11598\ : SRMux
    port map (
            O => \N__49473\,
            I => \N__49138\
        );

    \I__11597\ : SRMux
    port map (
            O => \N__49472\,
            I => \N__49138\
        );

    \I__11596\ : SRMux
    port map (
            O => \N__49471\,
            I => \N__49138\
        );

    \I__11595\ : SRMux
    port map (
            O => \N__49470\,
            I => \N__49138\
        );

    \I__11594\ : SRMux
    port map (
            O => \N__49469\,
            I => \N__49138\
        );

    \I__11593\ : SRMux
    port map (
            O => \N__49468\,
            I => \N__49138\
        );

    \I__11592\ : SRMux
    port map (
            O => \N__49467\,
            I => \N__49138\
        );

    \I__11591\ : SRMux
    port map (
            O => \N__49466\,
            I => \N__49138\
        );

    \I__11590\ : SRMux
    port map (
            O => \N__49465\,
            I => \N__49138\
        );

    \I__11589\ : SRMux
    port map (
            O => \N__49464\,
            I => \N__49138\
        );

    \I__11588\ : SRMux
    port map (
            O => \N__49463\,
            I => \N__49138\
        );

    \I__11587\ : SRMux
    port map (
            O => \N__49462\,
            I => \N__49138\
        );

    \I__11586\ : SRMux
    port map (
            O => \N__49461\,
            I => \N__49138\
        );

    \I__11585\ : SRMux
    port map (
            O => \N__49460\,
            I => \N__49138\
        );

    \I__11584\ : SRMux
    port map (
            O => \N__49459\,
            I => \N__49138\
        );

    \I__11583\ : SRMux
    port map (
            O => \N__49458\,
            I => \N__49138\
        );

    \I__11582\ : SRMux
    port map (
            O => \N__49457\,
            I => \N__49138\
        );

    \I__11581\ : SRMux
    port map (
            O => \N__49456\,
            I => \N__49138\
        );

    \I__11580\ : Glb2LocalMux
    port map (
            O => \N__49453\,
            I => \N__49138\
        );

    \I__11579\ : SRMux
    port map (
            O => \N__49452\,
            I => \N__49138\
        );

    \I__11578\ : SRMux
    port map (
            O => \N__49451\,
            I => \N__49138\
        );

    \I__11577\ : SRMux
    port map (
            O => \N__49450\,
            I => \N__49138\
        );

    \I__11576\ : SRMux
    port map (
            O => \N__49449\,
            I => \N__49138\
        );

    \I__11575\ : SRMux
    port map (
            O => \N__49448\,
            I => \N__49138\
        );

    \I__11574\ : Glb2LocalMux
    port map (
            O => \N__49445\,
            I => \N__49138\
        );

    \I__11573\ : SRMux
    port map (
            O => \N__49444\,
            I => \N__49138\
        );

    \I__11572\ : SRMux
    port map (
            O => \N__49443\,
            I => \N__49138\
        );

    \I__11571\ : SRMux
    port map (
            O => \N__49442\,
            I => \N__49138\
        );

    \I__11570\ : SRMux
    port map (
            O => \N__49441\,
            I => \N__49138\
        );

    \I__11569\ : SRMux
    port map (
            O => \N__49440\,
            I => \N__49138\
        );

    \I__11568\ : SRMux
    port map (
            O => \N__49439\,
            I => \N__49138\
        );

    \I__11567\ : SRMux
    port map (
            O => \N__49438\,
            I => \N__49138\
        );

    \I__11566\ : SRMux
    port map (
            O => \N__49437\,
            I => \N__49138\
        );

    \I__11565\ : SRMux
    port map (
            O => \N__49436\,
            I => \N__49138\
        );

    \I__11564\ : SRMux
    port map (
            O => \N__49435\,
            I => \N__49138\
        );

    \I__11563\ : SRMux
    port map (
            O => \N__49434\,
            I => \N__49138\
        );

    \I__11562\ : SRMux
    port map (
            O => \N__49433\,
            I => \N__49138\
        );

    \I__11561\ : SRMux
    port map (
            O => \N__49432\,
            I => \N__49138\
        );

    \I__11560\ : SRMux
    port map (
            O => \N__49431\,
            I => \N__49138\
        );

    \I__11559\ : SRMux
    port map (
            O => \N__49430\,
            I => \N__49138\
        );

    \I__11558\ : Glb2LocalMux
    port map (
            O => \N__49427\,
            I => \N__49138\
        );

    \I__11557\ : SRMux
    port map (
            O => \N__49426\,
            I => \N__49138\
        );

    \I__11556\ : SRMux
    port map (
            O => \N__49425\,
            I => \N__49138\
        );

    \I__11555\ : SRMux
    port map (
            O => \N__49424\,
            I => \N__49138\
        );

    \I__11554\ : SRMux
    port map (
            O => \N__49423\,
            I => \N__49138\
        );

    \I__11553\ : SRMux
    port map (
            O => \N__49422\,
            I => \N__49138\
        );

    \I__11552\ : SRMux
    port map (
            O => \N__49421\,
            I => \N__49138\
        );

    \I__11551\ : SRMux
    port map (
            O => \N__49420\,
            I => \N__49138\
        );

    \I__11550\ : Glb2LocalMux
    port map (
            O => \N__49417\,
            I => \N__49138\
        );

    \I__11549\ : SRMux
    port map (
            O => \N__49416\,
            I => \N__49138\
        );

    \I__11548\ : SRMux
    port map (
            O => \N__49415\,
            I => \N__49138\
        );

    \I__11547\ : SRMux
    port map (
            O => \N__49414\,
            I => \N__49138\
        );

    \I__11546\ : SRMux
    port map (
            O => \N__49413\,
            I => \N__49138\
        );

    \I__11545\ : SRMux
    port map (
            O => \N__49412\,
            I => \N__49138\
        );

    \I__11544\ : SRMux
    port map (
            O => \N__49411\,
            I => \N__49138\
        );

    \I__11543\ : SRMux
    port map (
            O => \N__49410\,
            I => \N__49138\
        );

    \I__11542\ : SRMux
    port map (
            O => \N__49409\,
            I => \N__49138\
        );

    \I__11541\ : SRMux
    port map (
            O => \N__49408\,
            I => \N__49138\
        );

    \I__11540\ : SRMux
    port map (
            O => \N__49407\,
            I => \N__49138\
        );

    \I__11539\ : SRMux
    port map (
            O => \N__49406\,
            I => \N__49138\
        );

    \I__11538\ : SRMux
    port map (
            O => \N__49405\,
            I => \N__49138\
        );

    \I__11537\ : GlobalMux
    port map (
            O => \N__49138\,
            I => \N__49135\
        );

    \I__11536\ : gio2CtrlBuf
    port map (
            O => \N__49135\,
            I => red_c_g
        );

    \I__11535\ : InMux
    port map (
            O => \N__49132\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__11534\ : InMux
    port map (
            O => \N__49129\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__11533\ : InMux
    port map (
            O => \N__49126\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__11532\ : CEMux
    port map (
            O => \N__49123\,
            I => \N__49117\
        );

    \I__11531\ : CEMux
    port map (
            O => \N__49122\,
            I => \N__49114\
        );

    \I__11530\ : CEMux
    port map (
            O => \N__49121\,
            I => \N__49111\
        );

    \I__11529\ : CEMux
    port map (
            O => \N__49120\,
            I => \N__49105\
        );

    \I__11528\ : LocalMux
    port map (
            O => \N__49117\,
            I => \N__49095\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__49114\,
            I => \N__49076\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__49111\,
            I => \N__49073\
        );

    \I__11525\ : CEMux
    port map (
            O => \N__49110\,
            I => \N__49070\
        );

    \I__11524\ : CEMux
    port map (
            O => \N__49109\,
            I => \N__49066\
        );

    \I__11523\ : CEMux
    port map (
            O => \N__49108\,
            I => \N__49063\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__49105\,
            I => \N__49060\
        );

    \I__11521\ : InMux
    port map (
            O => \N__49104\,
            I => \N__49051\
        );

    \I__11520\ : InMux
    port map (
            O => \N__49103\,
            I => \N__49051\
        );

    \I__11519\ : InMux
    port map (
            O => \N__49102\,
            I => \N__49051\
        );

    \I__11518\ : InMux
    port map (
            O => \N__49101\,
            I => \N__49051\
        );

    \I__11517\ : InMux
    port map (
            O => \N__49100\,
            I => \N__49044\
        );

    \I__11516\ : InMux
    port map (
            O => \N__49099\,
            I => \N__49044\
        );

    \I__11515\ : InMux
    port map (
            O => \N__49098\,
            I => \N__49044\
        );

    \I__11514\ : Span4Mux_h
    port map (
            O => \N__49095\,
            I => \N__49041\
        );

    \I__11513\ : InMux
    port map (
            O => \N__49094\,
            I => \N__49032\
        );

    \I__11512\ : InMux
    port map (
            O => \N__49093\,
            I => \N__49032\
        );

    \I__11511\ : InMux
    port map (
            O => \N__49092\,
            I => \N__49032\
        );

    \I__11510\ : InMux
    port map (
            O => \N__49091\,
            I => \N__49032\
        );

    \I__11509\ : InMux
    port map (
            O => \N__49090\,
            I => \N__49023\
        );

    \I__11508\ : InMux
    port map (
            O => \N__49089\,
            I => \N__49023\
        );

    \I__11507\ : InMux
    port map (
            O => \N__49088\,
            I => \N__49023\
        );

    \I__11506\ : InMux
    port map (
            O => \N__49087\,
            I => \N__49023\
        );

    \I__11505\ : InMux
    port map (
            O => \N__49086\,
            I => \N__49014\
        );

    \I__11504\ : InMux
    port map (
            O => \N__49085\,
            I => \N__49014\
        );

    \I__11503\ : InMux
    port map (
            O => \N__49084\,
            I => \N__49014\
        );

    \I__11502\ : InMux
    port map (
            O => \N__49083\,
            I => \N__49014\
        );

    \I__11501\ : InMux
    port map (
            O => \N__49082\,
            I => \N__49005\
        );

    \I__11500\ : InMux
    port map (
            O => \N__49081\,
            I => \N__49005\
        );

    \I__11499\ : InMux
    port map (
            O => \N__49080\,
            I => \N__49005\
        );

    \I__11498\ : InMux
    port map (
            O => \N__49079\,
            I => \N__49005\
        );

    \I__11497\ : Span4Mux_h
    port map (
            O => \N__49076\,
            I => \N__48998\
        );

    \I__11496\ : Span4Mux_h
    port map (
            O => \N__49073\,
            I => \N__48998\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__49070\,
            I => \N__48998\
        );

    \I__11494\ : CEMux
    port map (
            O => \N__49069\,
            I => \N__48995\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__49066\,
            I => \N__48990\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__49063\,
            I => \N__48987\
        );

    \I__11491\ : Span4Mux_v
    port map (
            O => \N__49060\,
            I => \N__48980\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__49051\,
            I => \N__48975\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__49044\,
            I => \N__48975\
        );

    \I__11488\ : Span4Mux_h
    port map (
            O => \N__49041\,
            I => \N__48964\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__49032\,
            I => \N__48964\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__49023\,
            I => \N__48964\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__49014\,
            I => \N__48964\
        );

    \I__11484\ : LocalMux
    port map (
            O => \N__49005\,
            I => \N__48964\
        );

    \I__11483\ : Span4Mux_v
    port map (
            O => \N__48998\,
            I => \N__48958\
        );

    \I__11482\ : LocalMux
    port map (
            O => \N__48995\,
            I => \N__48955\
        );

    \I__11481\ : InMux
    port map (
            O => \N__48994\,
            I => \N__48952\
        );

    \I__11480\ : CEMux
    port map (
            O => \N__48993\,
            I => \N__48948\
        );

    \I__11479\ : Span12Mux_h
    port map (
            O => \N__48990\,
            I => \N__48943\
        );

    \I__11478\ : Sp12to4
    port map (
            O => \N__48987\,
            I => \N__48943\
        );

    \I__11477\ : InMux
    port map (
            O => \N__48986\,
            I => \N__48934\
        );

    \I__11476\ : InMux
    port map (
            O => \N__48985\,
            I => \N__48934\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48984\,
            I => \N__48934\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48983\,
            I => \N__48934\
        );

    \I__11473\ : Span4Mux_h
    port map (
            O => \N__48980\,
            I => \N__48929\
        );

    \I__11472\ : Span4Mux_v
    port map (
            O => \N__48975\,
            I => \N__48929\
        );

    \I__11471\ : Span4Mux_v
    port map (
            O => \N__48964\,
            I => \N__48926\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48963\,
            I => \N__48919\
        );

    \I__11469\ : InMux
    port map (
            O => \N__48962\,
            I => \N__48919\
        );

    \I__11468\ : InMux
    port map (
            O => \N__48961\,
            I => \N__48919\
        );

    \I__11467\ : Span4Mux_h
    port map (
            O => \N__48958\,
            I => \N__48912\
        );

    \I__11466\ : Span4Mux_v
    port map (
            O => \N__48955\,
            I => \N__48912\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__48952\,
            I => \N__48912\
        );

    \I__11464\ : CEMux
    port map (
            O => \N__48951\,
            I => \N__48909\
        );

    \I__11463\ : LocalMux
    port map (
            O => \N__48948\,
            I => \N__48896\
        );

    \I__11462\ : Span12Mux_v
    port map (
            O => \N__48943\,
            I => \N__48896\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__48934\,
            I => \N__48896\
        );

    \I__11460\ : Sp12to4
    port map (
            O => \N__48929\,
            I => \N__48896\
        );

    \I__11459\ : Sp12to4
    port map (
            O => \N__48926\,
            I => \N__48896\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__48919\,
            I => \N__48896\
        );

    \I__11457\ : Span4Mux_v
    port map (
            O => \N__48912\,
            I => \N__48893\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__48909\,
            I => \N__48888\
        );

    \I__11455\ : Span12Mux_s9_h
    port map (
            O => \N__48896\,
            I => \N__48888\
        );

    \I__11454\ : Odrv4
    port map (
            O => \N__48893\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__11453\ : Odrv12
    port map (
            O => \N__48888\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__11452\ : InMux
    port map (
            O => \N__48883\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48880\,
            I => \N__48877\
        );

    \I__11450\ : LocalMux
    port map (
            O => \N__48877\,
            I => \N__48873\
        );

    \I__11449\ : InMux
    port map (
            O => \N__48876\,
            I => \N__48870\
        );

    \I__11448\ : Span4Mux_v
    port map (
            O => \N__48873\,
            I => \N__48867\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__48870\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__11446\ : Odrv4
    port map (
            O => \N__48867\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__11445\ : InMux
    port map (
            O => \N__48862\,
            I => \N__48858\
        );

    \I__11444\ : InMux
    port map (
            O => \N__48861\,
            I => \N__48855\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__48858\,
            I => \N__48852\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__48855\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__11441\ : Odrv12
    port map (
            O => \N__48852\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__11440\ : InMux
    port map (
            O => \N__48847\,
            I => \N__48844\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__48844\,
            I => \N__48841\
        );

    \I__11438\ : Span4Mux_h
    port map (
            O => \N__48841\,
            I => \N__48838\
        );

    \I__11437\ : Span4Mux_v
    port map (
            O => \N__48838\,
            I => \N__48835\
        );

    \I__11436\ : Odrv4
    port map (
            O => \N__48835\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df20\
        );

    \I__11435\ : InMux
    port map (
            O => \N__48832\,
            I => \N__48828\
        );

    \I__11434\ : InMux
    port map (
            O => \N__48831\,
            I => \N__48825\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__48828\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__48825\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__11431\ : InMux
    port map (
            O => \N__48820\,
            I => \N__48816\
        );

    \I__11430\ : InMux
    port map (
            O => \N__48819\,
            I => \N__48813\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__48816\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__48813\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__11427\ : InMux
    port map (
            O => \N__48808\,
            I => \N__48805\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__48805\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df26\
        );

    \I__11425\ : InMux
    port map (
            O => \N__48802\,
            I => \N__48798\
        );

    \I__11424\ : InMux
    port map (
            O => \N__48801\,
            I => \N__48795\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__48798\,
            I => \N__48792\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__48795\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__11421\ : Odrv4
    port map (
            O => \N__48792\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__11420\ : InMux
    port map (
            O => \N__48787\,
            I => \N__48783\
        );

    \I__11419\ : InMux
    port map (
            O => \N__48786\,
            I => \N__48780\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__48783\,
            I => \N__48777\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__48780\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__11416\ : Odrv4
    port map (
            O => \N__48777\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__11415\ : InMux
    port map (
            O => \N__48772\,
            I => \N__48769\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__48769\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df22\
        );

    \I__11413\ : InMux
    port map (
            O => \N__48766\,
            I => \N__48762\
        );

    \I__11412\ : InMux
    port map (
            O => \N__48765\,
            I => \N__48759\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__48762\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__48759\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__11409\ : InMux
    port map (
            O => \N__48754\,
            I => \N__48750\
        );

    \I__11408\ : InMux
    port map (
            O => \N__48753\,
            I => \N__48747\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__48750\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__48747\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__11405\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48739\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48739\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df28\
        );

    \I__11403\ : InMux
    port map (
            O => \N__48736\,
            I => \N__48731\
        );

    \I__11402\ : InMux
    port map (
            O => \N__48735\,
            I => \N__48728\
        );

    \I__11401\ : InMux
    port map (
            O => \N__48734\,
            I => \N__48725\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__48731\,
            I => \N__48722\
        );

    \I__11399\ : LocalMux
    port map (
            O => \N__48728\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__48725\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__11397\ : Odrv4
    port map (
            O => \N__48722\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__11396\ : CascadeMux
    port map (
            O => \N__48715\,
            I => \N__48712\
        );

    \I__11395\ : InMux
    port map (
            O => \N__48712\,
            I => \N__48707\
        );

    \I__11394\ : CascadeMux
    port map (
            O => \N__48711\,
            I => \N__48703\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48710\,
            I => \N__48700\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__48707\,
            I => \N__48697\
        );

    \I__11391\ : InMux
    port map (
            O => \N__48706\,
            I => \N__48694\
        );

    \I__11390\ : InMux
    port map (
            O => \N__48703\,
            I => \N__48691\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__48700\,
            I => \N__48686\
        );

    \I__11388\ : Span4Mux_h
    port map (
            O => \N__48697\,
            I => \N__48686\
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__48694\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__11386\ : LocalMux
    port map (
            O => \N__48691\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__11385\ : Odrv4
    port map (
            O => \N__48686\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__11384\ : InMux
    port map (
            O => \N__48679\,
            I => \N__48676\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__48676\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__11382\ : CascadeMux
    port map (
            O => \N__48673\,
            I => \N__48670\
        );

    \I__11381\ : InMux
    port map (
            O => \N__48670\,
            I => \N__48666\
        );

    \I__11380\ : InMux
    port map (
            O => \N__48669\,
            I => \N__48662\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__48666\,
            I => \N__48659\
        );

    \I__11378\ : InMux
    port map (
            O => \N__48665\,
            I => \N__48656\
        );

    \I__11377\ : LocalMux
    port map (
            O => \N__48662\,
            I => \N__48651\
        );

    \I__11376\ : Span4Mux_v
    port map (
            O => \N__48659\,
            I => \N__48651\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__48656\,
            I => \N__48648\
        );

    \I__11374\ : Odrv4
    port map (
            O => \N__48651\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__11373\ : Odrv4
    port map (
            O => \N__48648\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__11372\ : InMux
    port map (
            O => \N__48643\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__11371\ : InMux
    port map (
            O => \N__48640\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__11370\ : InMux
    port map (
            O => \N__48637\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__11369\ : InMux
    port map (
            O => \N__48634\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__11368\ : InMux
    port map (
            O => \N__48631\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__11367\ : InMux
    port map (
            O => \N__48628\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__11366\ : InMux
    port map (
            O => \N__48625\,
            I => \bfn_18_20_0_\
        );

    \I__11365\ : InMux
    port map (
            O => \N__48622\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__11364\ : InMux
    port map (
            O => \N__48619\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__11363\ : InMux
    port map (
            O => \N__48616\,
            I => \N__48612\
        );

    \I__11362\ : InMux
    port map (
            O => \N__48615\,
            I => \N__48609\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__48612\,
            I => \N__48606\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__48609\,
            I => \N__48601\
        );

    \I__11359\ : Span4Mux_v
    port map (
            O => \N__48606\,
            I => \N__48601\
        );

    \I__11358\ : Odrv4
    port map (
            O => \N__48601\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__11357\ : InMux
    port map (
            O => \N__48598\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__11356\ : InMux
    port map (
            O => \N__48595\,
            I => \N__48591\
        );

    \I__11355\ : InMux
    port map (
            O => \N__48594\,
            I => \N__48588\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__48591\,
            I => \N__48585\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__48588\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__11352\ : Odrv4
    port map (
            O => \N__48585\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__11351\ : InMux
    port map (
            O => \N__48580\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__11350\ : InMux
    port map (
            O => \N__48577\,
            I => \N__48573\
        );

    \I__11349\ : InMux
    port map (
            O => \N__48576\,
            I => \N__48570\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__48573\,
            I => \N__48567\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__48570\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__11346\ : Odrv4
    port map (
            O => \N__48567\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__11345\ : InMux
    port map (
            O => \N__48562\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__11344\ : InMux
    port map (
            O => \N__48559\,
            I => \N__48555\
        );

    \I__11343\ : InMux
    port map (
            O => \N__48558\,
            I => \N__48552\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__48555\,
            I => \N__48549\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__48552\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__11340\ : Odrv4
    port map (
            O => \N__48549\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__11339\ : InMux
    port map (
            O => \N__48544\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__11338\ : InMux
    port map (
            O => \N__48541\,
            I => \N__48537\
        );

    \I__11337\ : InMux
    port map (
            O => \N__48540\,
            I => \N__48534\
        );

    \I__11336\ : LocalMux
    port map (
            O => \N__48537\,
            I => \N__48531\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__48534\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__11334\ : Odrv4
    port map (
            O => \N__48531\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__11333\ : InMux
    port map (
            O => \N__48526\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__11332\ : CascadeMux
    port map (
            O => \N__48523\,
            I => \N__48520\
        );

    \I__11331\ : InMux
    port map (
            O => \N__48520\,
            I => \N__48514\
        );

    \I__11330\ : InMux
    port map (
            O => \N__48519\,
            I => \N__48514\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__48514\,
            I => \N__48510\
        );

    \I__11328\ : InMux
    port map (
            O => \N__48513\,
            I => \N__48507\
        );

    \I__11327\ : Span4Mux_h
    port map (
            O => \N__48510\,
            I => \N__48504\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__48507\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__11325\ : Odrv4
    port map (
            O => \N__48504\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__11324\ : InMux
    port map (
            O => \N__48499\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__11323\ : InMux
    port map (
            O => \N__48496\,
            I => \N__48489\
        );

    \I__11322\ : InMux
    port map (
            O => \N__48495\,
            I => \N__48489\
        );

    \I__11321\ : InMux
    port map (
            O => \N__48494\,
            I => \N__48486\
        );

    \I__11320\ : LocalMux
    port map (
            O => \N__48489\,
            I => \N__48483\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__48486\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__11318\ : Odrv4
    port map (
            O => \N__48483\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__11317\ : InMux
    port map (
            O => \N__48478\,
            I => \bfn_18_19_0_\
        );

    \I__11316\ : CascadeMux
    port map (
            O => \N__48475\,
            I => \N__48471\
        );

    \I__11315\ : InMux
    port map (
            O => \N__48474\,
            I => \N__48468\
        );

    \I__11314\ : InMux
    port map (
            O => \N__48471\,
            I => \N__48464\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__48468\,
            I => \N__48461\
        );

    \I__11312\ : InMux
    port map (
            O => \N__48467\,
            I => \N__48458\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__48464\,
            I => \N__48455\
        );

    \I__11310\ : Span4Mux_h
    port map (
            O => \N__48461\,
            I => \N__48452\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__48458\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__11308\ : Odrv12
    port map (
            O => \N__48455\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__11307\ : Odrv4
    port map (
            O => \N__48452\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__11306\ : InMux
    port map (
            O => \N__48445\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__11305\ : InMux
    port map (
            O => \N__48442\,
            I => \N__48439\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__48439\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28\
        );

    \I__11303\ : CascadeMux
    port map (
            O => \N__48436\,
            I => \N__48432\
        );

    \I__11302\ : InMux
    port map (
            O => \N__48435\,
            I => \N__48429\
        );

    \I__11301\ : InMux
    port map (
            O => \N__48432\,
            I => \N__48426\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__48429\,
            I => \N__48423\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__48426\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__11298\ : Odrv4
    port map (
            O => \N__48423\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__11297\ : InMux
    port map (
            O => \N__48418\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__11296\ : InMux
    port map (
            O => \N__48415\,
            I => \N__48411\
        );

    \I__11295\ : InMux
    port map (
            O => \N__48414\,
            I => \N__48408\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__48411\,
            I => \N__48405\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__48408\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__11292\ : Odrv4
    port map (
            O => \N__48405\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__11291\ : InMux
    port map (
            O => \N__48400\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__11290\ : InMux
    port map (
            O => \N__48397\,
            I => \N__48393\
        );

    \I__11289\ : InMux
    port map (
            O => \N__48396\,
            I => \N__48390\
        );

    \I__11288\ : LocalMux
    port map (
            O => \N__48393\,
            I => \N__48387\
        );

    \I__11287\ : LocalMux
    port map (
            O => \N__48390\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__11286\ : Odrv4
    port map (
            O => \N__48387\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__11285\ : InMux
    port map (
            O => \N__48382\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__11284\ : InMux
    port map (
            O => \N__48379\,
            I => \N__48375\
        );

    \I__11283\ : InMux
    port map (
            O => \N__48378\,
            I => \N__48372\
        );

    \I__11282\ : LocalMux
    port map (
            O => \N__48375\,
            I => \N__48369\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__48372\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__11280\ : Odrv4
    port map (
            O => \N__48369\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__11279\ : InMux
    port map (
            O => \N__48364\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__11278\ : InMux
    port map (
            O => \N__48361\,
            I => \N__48357\
        );

    \I__11277\ : InMux
    port map (
            O => \N__48360\,
            I => \N__48354\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__48357\,
            I => \N__48351\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__48354\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__11274\ : Odrv4
    port map (
            O => \N__48351\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__11273\ : InMux
    port map (
            O => \N__48346\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__11272\ : InMux
    port map (
            O => \N__48343\,
            I => \N__48339\
        );

    \I__11271\ : InMux
    port map (
            O => \N__48342\,
            I => \N__48336\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__48339\,
            I => \N__48333\
        );

    \I__11269\ : LocalMux
    port map (
            O => \N__48336\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__11268\ : Odrv4
    port map (
            O => \N__48333\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__11267\ : InMux
    port map (
            O => \N__48328\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__11266\ : InMux
    port map (
            O => \N__48325\,
            I => \N__48321\
        );

    \I__11265\ : InMux
    port map (
            O => \N__48324\,
            I => \N__48318\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__48321\,
            I => \N__48315\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__48318\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__11262\ : Odrv4
    port map (
            O => \N__48315\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__11261\ : InMux
    port map (
            O => \N__48310\,
            I => \bfn_18_18_0_\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48307\,
            I => \N__48304\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__48304\,
            I => \N__48300\
        );

    \I__11258\ : InMux
    port map (
            O => \N__48303\,
            I => \N__48297\
        );

    \I__11257\ : Span4Mux_v
    port map (
            O => \N__48300\,
            I => \N__48294\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__48297\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__11255\ : Odrv4
    port map (
            O => \N__48294\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__11254\ : InMux
    port map (
            O => \N__48289\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__11253\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48283\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__48283\,
            I => \N__48280\
        );

    \I__11251\ : Span4Mux_v
    port map (
            O => \N__48280\,
            I => \N__48276\
        );

    \I__11250\ : InMux
    port map (
            O => \N__48279\,
            I => \N__48273\
        );

    \I__11249\ : Span4Mux_h
    port map (
            O => \N__48276\,
            I => \N__48270\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__48273\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__11247\ : Odrv4
    port map (
            O => \N__48270\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__11246\ : InMux
    port map (
            O => \N__48265\,
            I => \bfn_18_16_0_\
        );

    \I__11245\ : InMux
    port map (
            O => \N__48262\,
            I => \N__48258\
        );

    \I__11244\ : InMux
    port map (
            O => \N__48261\,
            I => \N__48255\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__48258\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__48255\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__11241\ : InMux
    port map (
            O => \N__48250\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__11240\ : InMux
    port map (
            O => \N__48247\,
            I => \N__48243\
        );

    \I__11239\ : InMux
    port map (
            O => \N__48246\,
            I => \N__48240\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__48243\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__48240\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__11236\ : InMux
    port map (
            O => \N__48235\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__11235\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48228\
        );

    \I__11234\ : InMux
    port map (
            O => \N__48231\,
            I => \N__48225\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__48228\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__48225\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__11231\ : InMux
    port map (
            O => \N__48220\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__11230\ : InMux
    port map (
            O => \N__48217\,
            I => \N__48213\
        );

    \I__11229\ : InMux
    port map (
            O => \N__48216\,
            I => \N__48210\
        );

    \I__11228\ : LocalMux
    port map (
            O => \N__48213\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__48210\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__11226\ : InMux
    port map (
            O => \N__48205\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__11225\ : InMux
    port map (
            O => \N__48202\,
            I => \N__48197\
        );

    \I__11224\ : InMux
    port map (
            O => \N__48201\,
            I => \N__48194\
        );

    \I__11223\ : InMux
    port map (
            O => \N__48200\,
            I => \N__48191\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__48197\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__48194\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__48191\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__11219\ : InMux
    port map (
            O => \N__48184\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__11218\ : InMux
    port map (
            O => \N__48181\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__11217\ : CascadeMux
    port map (
            O => \N__48178\,
            I => \N__48175\
        );

    \I__11216\ : InMux
    port map (
            O => \N__48175\,
            I => \N__48172\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__48172\,
            I => \N__48167\
        );

    \I__11214\ : CascadeMux
    port map (
            O => \N__48171\,
            I => \N__48163\
        );

    \I__11213\ : InMux
    port map (
            O => \N__48170\,
            I => \N__48160\
        );

    \I__11212\ : Span4Mux_h
    port map (
            O => \N__48167\,
            I => \N__48157\
        );

    \I__11211\ : InMux
    port map (
            O => \N__48166\,
            I => \N__48154\
        );

    \I__11210\ : InMux
    port map (
            O => \N__48163\,
            I => \N__48151\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__48160\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__11208\ : Odrv4
    port map (
            O => \N__48157\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__48154\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__48151\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__11205\ : InMux
    port map (
            O => \N__48142\,
            I => \N__48137\
        );

    \I__11204\ : InMux
    port map (
            O => \N__48141\,
            I => \N__48134\
        );

    \I__11203\ : InMux
    port map (
            O => \N__48140\,
            I => \N__48131\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__48137\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__48134\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__48131\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__11199\ : CascadeMux
    port map (
            O => \N__48124\,
            I => \N__48121\
        );

    \I__11198\ : InMux
    port map (
            O => \N__48121\,
            I => \N__48118\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__48118\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__11196\ : InMux
    port map (
            O => \N__48115\,
            I => \N__48111\
        );

    \I__11195\ : InMux
    port map (
            O => \N__48114\,
            I => \N__48108\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__48111\,
            I => \N__48105\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__48108\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__11192\ : Odrv4
    port map (
            O => \N__48105\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__11191\ : InMux
    port map (
            O => \N__48100\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__11190\ : CascadeMux
    port map (
            O => \N__48097\,
            I => \N__48094\
        );

    \I__11189\ : InMux
    port map (
            O => \N__48094\,
            I => \N__48088\
        );

    \I__11188\ : InMux
    port map (
            O => \N__48093\,
            I => \N__48088\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__48088\,
            I => \N__48084\
        );

    \I__11186\ : InMux
    port map (
            O => \N__48087\,
            I => \N__48081\
        );

    \I__11185\ : Span4Mux_v
    port map (
            O => \N__48084\,
            I => \N__48078\
        );

    \I__11184\ : LocalMux
    port map (
            O => \N__48081\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__11183\ : Odrv4
    port map (
            O => \N__48078\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__11182\ : InMux
    port map (
            O => \N__48073\,
            I => \bfn_18_15_0_\
        );

    \I__11181\ : InMux
    port map (
            O => \N__48070\,
            I => \N__48064\
        );

    \I__11180\ : InMux
    port map (
            O => \N__48069\,
            I => \N__48064\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__48064\,
            I => \N__48060\
        );

    \I__11178\ : InMux
    port map (
            O => \N__48063\,
            I => \N__48057\
        );

    \I__11177\ : Span4Mux_v
    port map (
            O => \N__48060\,
            I => \N__48054\
        );

    \I__11176\ : LocalMux
    port map (
            O => \N__48057\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__11175\ : Odrv4
    port map (
            O => \N__48054\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__11174\ : InMux
    port map (
            O => \N__48049\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__11173\ : CascadeMux
    port map (
            O => \N__48046\,
            I => \N__48043\
        );

    \I__11172\ : InMux
    port map (
            O => \N__48043\,
            I => \N__48037\
        );

    \I__11171\ : InMux
    port map (
            O => \N__48042\,
            I => \N__48037\
        );

    \I__11170\ : LocalMux
    port map (
            O => \N__48037\,
            I => \N__48033\
        );

    \I__11169\ : InMux
    port map (
            O => \N__48036\,
            I => \N__48030\
        );

    \I__11168\ : Span4Mux_h
    port map (
            O => \N__48033\,
            I => \N__48027\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__48030\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__11166\ : Odrv4
    port map (
            O => \N__48027\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__11165\ : InMux
    port map (
            O => \N__48022\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__11164\ : InMux
    port map (
            O => \N__48019\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__11163\ : InMux
    port map (
            O => \N__48016\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__11162\ : InMux
    port map (
            O => \N__48013\,
            I => \N__48010\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__48010\,
            I => \N__48006\
        );

    \I__11160\ : InMux
    port map (
            O => \N__48009\,
            I => \N__48003\
        );

    \I__11159\ : Span4Mux_v
    port map (
            O => \N__48006\,
            I => \N__48000\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__48003\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__11157\ : Odrv4
    port map (
            O => \N__48000\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__11156\ : InMux
    port map (
            O => \N__47995\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__11155\ : InMux
    port map (
            O => \N__47992\,
            I => \N__47989\
        );

    \I__11154\ : LocalMux
    port map (
            O => \N__47989\,
            I => \N__47986\
        );

    \I__11153\ : Span4Mux_v
    port map (
            O => \N__47986\,
            I => \N__47982\
        );

    \I__11152\ : InMux
    port map (
            O => \N__47985\,
            I => \N__47979\
        );

    \I__11151\ : Span4Mux_h
    port map (
            O => \N__47982\,
            I => \N__47976\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__47979\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__11149\ : Odrv4
    port map (
            O => \N__47976\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__11148\ : InMux
    port map (
            O => \N__47971\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__11147\ : InMux
    port map (
            O => \N__47968\,
            I => \N__47965\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__47965\,
            I => \N__47962\
        );

    \I__11145\ : Span4Mux_h
    port map (
            O => \N__47962\,
            I => \N__47958\
        );

    \I__11144\ : InMux
    port map (
            O => \N__47961\,
            I => \N__47955\
        );

    \I__11143\ : Span4Mux_v
    port map (
            O => \N__47958\,
            I => \N__47952\
        );

    \I__11142\ : LocalMux
    port map (
            O => \N__47955\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__11141\ : Odrv4
    port map (
            O => \N__47952\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__11140\ : InMux
    port map (
            O => \N__47947\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__11139\ : InMux
    port map (
            O => \N__47944\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__11138\ : InMux
    port map (
            O => \N__47941\,
            I => \N__47937\
        );

    \I__11137\ : InMux
    port map (
            O => \N__47940\,
            I => \N__47934\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__47937\,
            I => \N__47931\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__47934\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__11134\ : Odrv12
    port map (
            O => \N__47931\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47926\,
            I => \bfn_18_14_0_\
        );

    \I__11132\ : InMux
    port map (
            O => \N__47923\,
            I => \N__47919\
        );

    \I__11131\ : InMux
    port map (
            O => \N__47922\,
            I => \N__47916\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__47919\,
            I => \N__47913\
        );

    \I__11129\ : LocalMux
    port map (
            O => \N__47916\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__11128\ : Odrv12
    port map (
            O => \N__47913\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__11127\ : InMux
    port map (
            O => \N__47908\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__11126\ : InMux
    port map (
            O => \N__47905\,
            I => \N__47901\
        );

    \I__11125\ : InMux
    port map (
            O => \N__47904\,
            I => \N__47898\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__47901\,
            I => \N__47895\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__47898\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__11122\ : Odrv4
    port map (
            O => \N__47895\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__11121\ : InMux
    port map (
            O => \N__47890\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__11120\ : InMux
    port map (
            O => \N__47887\,
            I => \N__47883\
        );

    \I__11119\ : InMux
    port map (
            O => \N__47886\,
            I => \N__47880\
        );

    \I__11118\ : LocalMux
    port map (
            O => \N__47883\,
            I => \N__47877\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__47880\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__11116\ : Odrv4
    port map (
            O => \N__47877\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__11115\ : InMux
    port map (
            O => \N__47872\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__11114\ : InMux
    port map (
            O => \N__47869\,
            I => \N__47865\
        );

    \I__11113\ : InMux
    port map (
            O => \N__47868\,
            I => \N__47862\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__47865\,
            I => \N__47859\
        );

    \I__11111\ : LocalMux
    port map (
            O => \N__47862\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__11110\ : Odrv4
    port map (
            O => \N__47859\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__11109\ : InMux
    port map (
            O => \N__47854\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47851\,
            I => \N__47847\
        );

    \I__11107\ : InMux
    port map (
            O => \N__47850\,
            I => \N__47844\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__47847\,
            I => \N__47841\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__47844\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__11104\ : Odrv4
    port map (
            O => \N__47841\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__11103\ : InMux
    port map (
            O => \N__47836\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__11102\ : InMux
    port map (
            O => \N__47833\,
            I => \N__47829\
        );

    \I__11101\ : InMux
    port map (
            O => \N__47832\,
            I => \N__47826\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__47829\,
            I => \N__47823\
        );

    \I__11099\ : LocalMux
    port map (
            O => \N__47826\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__11098\ : Odrv12
    port map (
            O => \N__47823\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__11097\ : InMux
    port map (
            O => \N__47818\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__11096\ : InMux
    port map (
            O => \N__47815\,
            I => \N__47808\
        );

    \I__11095\ : InMux
    port map (
            O => \N__47814\,
            I => \N__47808\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47813\,
            I => \N__47805\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__47808\,
            I => \N__47802\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__47805\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__11091\ : Odrv4
    port map (
            O => \N__47802\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__11090\ : InMux
    port map (
            O => \N__47797\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__11089\ : InMux
    port map (
            O => \N__47794\,
            I => \N__47786\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47793\,
            I => \N__47786\
        );

    \I__11087\ : InMux
    port map (
            O => \N__47792\,
            I => \N__47781\
        );

    \I__11086\ : InMux
    port map (
            O => \N__47791\,
            I => \N__47781\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47786\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__47781\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\
        );

    \I__11083\ : CascadeMux
    port map (
            O => \N__47776\,
            I => \N__47772\
        );

    \I__11082\ : InMux
    port map (
            O => \N__47775\,
            I => \N__47767\
        );

    \I__11081\ : InMux
    port map (
            O => \N__47772\,
            I => \N__47767\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__47767\,
            I => \N__47764\
        );

    \I__11079\ : Span4Mux_h
    port map (
            O => \N__47764\,
            I => \N__47759\
        );

    \I__11078\ : InMux
    port map (
            O => \N__47763\,
            I => \N__47756\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47762\,
            I => \N__47753\
        );

    \I__11076\ : Odrv4
    port map (
            O => \N__47759\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__47756\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__47753\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\
        );

    \I__11073\ : CascadeMux
    port map (
            O => \N__47746\,
            I => \delay_measurement_inst.delay_tr_timer.N_362_cascade_\
        );

    \I__11072\ : InMux
    port map (
            O => \N__47743\,
            I => \N__47739\
        );

    \I__11071\ : CascadeMux
    port map (
            O => \N__47742\,
            I => \N__47735\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__47739\,
            I => \N__47731\
        );

    \I__11069\ : InMux
    port map (
            O => \N__47738\,
            I => \N__47724\
        );

    \I__11068\ : InMux
    port map (
            O => \N__47735\,
            I => \N__47724\
        );

    \I__11067\ : InMux
    port map (
            O => \N__47734\,
            I => \N__47724\
        );

    \I__11066\ : Odrv4
    port map (
            O => \N__47731\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__47724\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\
        );

    \I__11064\ : InMux
    port map (
            O => \N__47719\,
            I => \N__47715\
        );

    \I__11063\ : InMux
    port map (
            O => \N__47718\,
            I => \N__47712\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__47715\,
            I => \N__47708\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__47712\,
            I => \N__47705\
        );

    \I__11060\ : InMux
    port map (
            O => \N__47711\,
            I => \N__47702\
        );

    \I__11059\ : Span4Mux_v
    port map (
            O => \N__47708\,
            I => \N__47697\
        );

    \I__11058\ : Span4Mux_v
    port map (
            O => \N__47705\,
            I => \N__47697\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__47702\,
            I => \N__47694\
        );

    \I__11056\ : Odrv4
    port map (
            O => \N__47697\,
            I => \delay_measurement_inst.N_365\
        );

    \I__11055\ : Odrv4
    port map (
            O => \N__47694\,
            I => \delay_measurement_inst.N_365\
        );

    \I__11054\ : InMux
    port map (
            O => \N__47689\,
            I => \N__47686\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__47686\,
            I => \N__47683\
        );

    \I__11052\ : Odrv4
    port map (
            O => \N__47683\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__11051\ : CascadeMux
    port map (
            O => \N__47680\,
            I => \N__47676\
        );

    \I__11050\ : InMux
    port map (
            O => \N__47679\,
            I => \N__47673\
        );

    \I__11049\ : InMux
    port map (
            O => \N__47676\,
            I => \N__47670\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__47673\,
            I => \N__47664\
        );

    \I__11047\ : LocalMux
    port map (
            O => \N__47670\,
            I => \N__47664\
        );

    \I__11046\ : InMux
    port map (
            O => \N__47669\,
            I => \N__47661\
        );

    \I__11045\ : Odrv4
    port map (
            O => \N__47664\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__47661\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__11043\ : InMux
    port map (
            O => \N__47656\,
            I => \N__47652\
        );

    \I__11042\ : InMux
    port map (
            O => \N__47655\,
            I => \N__47649\
        );

    \I__11041\ : LocalMux
    port map (
            O => \N__47652\,
            I => \N__47646\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__47649\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__11039\ : Odrv12
    port map (
            O => \N__47646\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__11038\ : InMux
    port map (
            O => \N__47641\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__11037\ : CascadeMux
    port map (
            O => \N__47638\,
            I => \N__47635\
        );

    \I__11036\ : InMux
    port map (
            O => \N__47635\,
            I => \N__47632\
        );

    \I__11035\ : LocalMux
    port map (
            O => \N__47632\,
            I => \N__47629\
        );

    \I__11034\ : Span4Mux_h
    port map (
            O => \N__47629\,
            I => \N__47626\
        );

    \I__11033\ : Odrv4
    port map (
            O => \N__47626\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28\
        );

    \I__11032\ : InMux
    port map (
            O => \N__47623\,
            I => \N__47619\
        );

    \I__11031\ : InMux
    port map (
            O => \N__47622\,
            I => \N__47616\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__47619\,
            I => \N__47613\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__47616\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__11028\ : Odrv4
    port map (
            O => \N__47613\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__11027\ : InMux
    port map (
            O => \N__47608\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__11026\ : InMux
    port map (
            O => \N__47605\,
            I => \N__47602\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__47602\,
            I => \N__47598\
        );

    \I__11024\ : InMux
    port map (
            O => \N__47601\,
            I => \N__47595\
        );

    \I__11023\ : Sp12to4
    port map (
            O => \N__47598\,
            I => \N__47592\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__47595\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__11021\ : Odrv12
    port map (
            O => \N__47592\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__11020\ : InMux
    port map (
            O => \N__47587\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__11019\ : InMux
    port map (
            O => \N__47584\,
            I => \N__47580\
        );

    \I__11018\ : InMux
    port map (
            O => \N__47583\,
            I => \N__47577\
        );

    \I__11017\ : LocalMux
    port map (
            O => \N__47580\,
            I => \N__47574\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__47577\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__11015\ : Odrv12
    port map (
            O => \N__47574\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__11014\ : InMux
    port map (
            O => \N__47569\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__11013\ : InMux
    port map (
            O => \N__47566\,
            I => \N__47562\
        );

    \I__11012\ : InMux
    port map (
            O => \N__47565\,
            I => \N__47559\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__47562\,
            I => \N__47556\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__47559\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__11009\ : Odrv4
    port map (
            O => \N__47556\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__11008\ : InMux
    port map (
            O => \N__47551\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__11007\ : InMux
    port map (
            O => \N__47548\,
            I => \N__47545\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__47545\,
            I => \N__47541\
        );

    \I__11005\ : InMux
    port map (
            O => \N__47544\,
            I => \N__47538\
        );

    \I__11004\ : Span4Mux_h
    port map (
            O => \N__47541\,
            I => \N__47535\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__47538\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__11002\ : Odrv4
    port map (
            O => \N__47535\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__11001\ : InMux
    port map (
            O => \N__47530\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__11000\ : InMux
    port map (
            O => \N__47527\,
            I => \N__47523\
        );

    \I__10999\ : InMux
    port map (
            O => \N__47526\,
            I => \N__47520\
        );

    \I__10998\ : LocalMux
    port map (
            O => \N__47523\,
            I => \N__47517\
        );

    \I__10997\ : LocalMux
    port map (
            O => \N__47520\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10996\ : Odrv12
    port map (
            O => \N__47517\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10995\ : CascadeMux
    port map (
            O => \N__47512\,
            I => \N__47508\
        );

    \I__10994\ : InMux
    port map (
            O => \N__47511\,
            I => \N__47505\
        );

    \I__10993\ : InMux
    port map (
            O => \N__47508\,
            I => \N__47502\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__47505\,
            I => \N__47499\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__47502\,
            I => \N__47495\
        );

    \I__10990\ : Span4Mux_v
    port map (
            O => \N__47499\,
            I => \N__47492\
        );

    \I__10989\ : InMux
    port map (
            O => \N__47498\,
            I => \N__47489\
        );

    \I__10988\ : Span4Mux_v
    port map (
            O => \N__47495\,
            I => \N__47486\
        );

    \I__10987\ : Odrv4
    port map (
            O => \N__47492\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__47489\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10985\ : Odrv4
    port map (
            O => \N__47486\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10984\ : CEMux
    port map (
            O => \N__47479\,
            I => \N__47464\
        );

    \I__10983\ : CEMux
    port map (
            O => \N__47478\,
            I => \N__47464\
        );

    \I__10982\ : CEMux
    port map (
            O => \N__47477\,
            I => \N__47464\
        );

    \I__10981\ : CEMux
    port map (
            O => \N__47476\,
            I => \N__47464\
        );

    \I__10980\ : CEMux
    port map (
            O => \N__47475\,
            I => \N__47464\
        );

    \I__10979\ : GlobalMux
    port map (
            O => \N__47464\,
            I => \N__47461\
        );

    \I__10978\ : gio2CtrlBuf
    port map (
            O => \N__47461\,
            I => \delay_measurement_inst.delay_tr_timer.N_399_i_g\
        );

    \I__10977\ : CascadeMux
    port map (
            O => \N__47458\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\
        );

    \I__10976\ : CascadeMux
    port map (
            O => \N__47455\,
            I => \N__47452\
        );

    \I__10975\ : InMux
    port map (
            O => \N__47452\,
            I => \N__47448\
        );

    \I__10974\ : InMux
    port map (
            O => \N__47451\,
            I => \N__47445\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__47448\,
            I => \N__47442\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__47445\,
            I => \N__47439\
        );

    \I__10971\ : Span4Mux_h
    port map (
            O => \N__47442\,
            I => \N__47436\
        );

    \I__10970\ : Span4Mux_h
    port map (
            O => \N__47439\,
            I => \N__47433\
        );

    \I__10969\ : Odrv4
    port map (
            O => \N__47436\,
            I => \delay_measurement_inst.delay_tr_timer.N_394\
        );

    \I__10968\ : Odrv4
    port map (
            O => \N__47433\,
            I => \delay_measurement_inst.delay_tr_timer.N_394\
        );

    \I__10967\ : InMux
    port map (
            O => \N__47428\,
            I => \N__47425\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__47425\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\
        );

    \I__10965\ : InMux
    port map (
            O => \N__47422\,
            I => \N__47418\
        );

    \I__10964\ : InMux
    port map (
            O => \N__47421\,
            I => \N__47415\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__47418\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__47415\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__10961\ : CascadeMux
    port map (
            O => \N__47410\,
            I => \N__47407\
        );

    \I__10960\ : InMux
    port map (
            O => \N__47407\,
            I => \N__47403\
        );

    \I__10959\ : InMux
    port map (
            O => \N__47406\,
            I => \N__47400\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__47403\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__47400\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__10956\ : InMux
    port map (
            O => \N__47395\,
            I => \N__47392\
        );

    \I__10955\ : LocalMux
    port map (
            O => \N__47392\,
            I => \N__47389\
        );

    \I__10954\ : Odrv4
    port map (
            O => \N__47389\,
            I => \delay_measurement_inst.delay_tr_timer.N_346\
        );

    \I__10953\ : CascadeMux
    port map (
            O => \N__47386\,
            I => \N__47383\
        );

    \I__10952\ : InMux
    port map (
            O => \N__47383\,
            I => \N__47378\
        );

    \I__10951\ : InMux
    port map (
            O => \N__47382\,
            I => \N__47373\
        );

    \I__10950\ : InMux
    port map (
            O => \N__47381\,
            I => \N__47373\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__47378\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__47373\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__10947\ : CascadeMux
    port map (
            O => \N__47368\,
            I => \N__47365\
        );

    \I__10946\ : InMux
    port map (
            O => \N__47365\,
            I => \N__47361\
        );

    \I__10945\ : CascadeMux
    port map (
            O => \N__47364\,
            I => \N__47358\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__47361\,
            I => \N__47355\
        );

    \I__10943\ : InMux
    port map (
            O => \N__47358\,
            I => \N__47352\
        );

    \I__10942\ : Span12Mux_h
    port map (
            O => \N__47355\,
            I => \N__47348\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__47352\,
            I => \N__47345\
        );

    \I__10940\ : InMux
    port map (
            O => \N__47351\,
            I => \N__47342\
        );

    \I__10939\ : Odrv12
    port map (
            O => \N__47348\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__10938\ : Odrv4
    port map (
            O => \N__47345\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__47342\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__10936\ : CascadeMux
    port map (
            O => \N__47335\,
            I => \delay_measurement_inst.delay_tr_timer.N_346_cascade_\
        );

    \I__10935\ : CascadeMux
    port map (
            O => \N__47332\,
            I => \N__47329\
        );

    \I__10934\ : InMux
    port map (
            O => \N__47329\,
            I => \N__47326\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__47326\,
            I => \N__47323\
        );

    \I__10932\ : Span4Mux_h
    port map (
            O => \N__47323\,
            I => \N__47319\
        );

    \I__10931\ : InMux
    port map (
            O => \N__47322\,
            I => \N__47316\
        );

    \I__10930\ : Odrv4
    port map (
            O => \N__47319\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__47316\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__10928\ : InMux
    port map (
            O => \N__47311\,
            I => \N__47308\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__47308\,
            I => \N__47305\
        );

    \I__10926\ : Odrv4
    port map (
            O => \N__47305\,
            I => \delay_measurement_inst.delay_tr_timer.N_349\
        );

    \I__10925\ : CascadeMux
    port map (
            O => \N__47302\,
            I => \N__47299\
        );

    \I__10924\ : InMux
    port map (
            O => \N__47299\,
            I => \N__47296\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__47296\,
            I => \N__47293\
        );

    \I__10922\ : Span4Mux_h
    port map (
            O => \N__47293\,
            I => \N__47288\
        );

    \I__10921\ : InMux
    port map (
            O => \N__47292\,
            I => \N__47285\
        );

    \I__10920\ : InMux
    port map (
            O => \N__47291\,
            I => \N__47282\
        );

    \I__10919\ : Odrv4
    port map (
            O => \N__47288\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__47285\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__47282\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__10916\ : InMux
    port map (
            O => \N__47275\,
            I => \N__47272\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__47272\,
            I => \N__47269\
        );

    \I__10914\ : Span4Mux_h
    port map (
            O => \N__47269\,
            I => \N__47266\
        );

    \I__10913\ : Span4Mux_h
    port map (
            O => \N__47266\,
            I => \N__47261\
        );

    \I__10912\ : InMux
    port map (
            O => \N__47265\,
            I => \N__47258\
        );

    \I__10911\ : InMux
    port map (
            O => \N__47264\,
            I => \N__47255\
        );

    \I__10910\ : Odrv4
    port map (
            O => \N__47261\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__47258\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__47255\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__10907\ : CascadeMux
    port map (
            O => \N__47248\,
            I => \delay_measurement_inst.delay_tr_timer.N_349_cascade_\
        );

    \I__10906\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47242\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__47242\,
            I => \N__47239\
        );

    \I__10904\ : Span4Mux_h
    port map (
            O => \N__47239\,
            I => \N__47236\
        );

    \I__10903\ : Odrv4
    port map (
            O => \N__47236\,
            I => \delay_measurement_inst.delay_tr_timer.N_351\
        );

    \I__10902\ : InMux
    port map (
            O => \N__47233\,
            I => \N__47230\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__47230\,
            I => \N__47227\
        );

    \I__10900\ : Span4Mux_v
    port map (
            O => \N__47227\,
            I => \N__47222\
        );

    \I__10899\ : InMux
    port map (
            O => \N__47226\,
            I => \N__47217\
        );

    \I__10898\ : InMux
    port map (
            O => \N__47225\,
            I => \N__47217\
        );

    \I__10897\ : Odrv4
    port map (
            O => \N__47222\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__47217\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__10895\ : InMux
    port map (
            O => \N__47212\,
            I => \N__47209\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__47209\,
            I => \N__47204\
        );

    \I__10893\ : InMux
    port map (
            O => \N__47208\,
            I => \N__47199\
        );

    \I__10892\ : InMux
    port map (
            O => \N__47207\,
            I => \N__47199\
        );

    \I__10891\ : Odrv4
    port map (
            O => \N__47204\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__47199\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__10889\ : CascadeMux
    port map (
            O => \N__47194\,
            I => \N__47190\
        );

    \I__10888\ : InMux
    port map (
            O => \N__47193\,
            I => \N__47186\
        );

    \I__10887\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47183\
        );

    \I__10886\ : InMux
    port map (
            O => \N__47189\,
            I => \N__47180\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__47186\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__47183\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__47180\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__10882\ : InMux
    port map (
            O => \N__47173\,
            I => \N__47168\
        );

    \I__10881\ : InMux
    port map (
            O => \N__47172\,
            I => \N__47163\
        );

    \I__10880\ : InMux
    port map (
            O => \N__47171\,
            I => \N__47163\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__47168\,
            I => \N__47160\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__47163\,
            I => \N__47157\
        );

    \I__10877\ : Odrv12
    port map (
            O => \N__47160\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10876\ : Odrv4
    port map (
            O => \N__47157\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10875\ : InMux
    port map (
            O => \N__47152\,
            I => \N__47149\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__47149\,
            I => \N__47146\
        );

    \I__10873\ : Span4Mux_h
    port map (
            O => \N__47146\,
            I => \N__47143\
        );

    \I__10872\ : Odrv4
    port map (
            O => \N__47143\,
            I => \delay_measurement_inst.delay_tr_timer.N_362\
        );

    \I__10871\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47137\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__47137\,
            I => \N__47134\
        );

    \I__10869\ : Odrv12
    port map (
            O => \N__47134\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__10868\ : InMux
    port map (
            O => \N__47131\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28\
        );

    \I__10867\ : InMux
    port map (
            O => \N__47128\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__10866\ : InMux
    port map (
            O => \N__47125\,
            I => \N__47119\
        );

    \I__10865\ : InMux
    port map (
            O => \N__47124\,
            I => \N__47119\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__47119\,
            I => \N__47116\
        );

    \I__10863\ : Odrv12
    port map (
            O => \N__47116\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__10862\ : InMux
    port map (
            O => \N__47113\,
            I => \N__47108\
        );

    \I__10861\ : InMux
    port map (
            O => \N__47112\,
            I => \N__47102\
        );

    \I__10860\ : InMux
    port map (
            O => \N__47111\,
            I => \N__47099\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__47108\,
            I => \N__47094\
        );

    \I__10858\ : InMux
    port map (
            O => \N__47107\,
            I => \N__47089\
        );

    \I__10857\ : InMux
    port map (
            O => \N__47106\,
            I => \N__47089\
        );

    \I__10856\ : CascadeMux
    port map (
            O => \N__47105\,
            I => \N__47080\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__47102\,
            I => \N__47073\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__47099\,
            I => \N__47052\
        );

    \I__10853\ : InMux
    port map (
            O => \N__47098\,
            I => \N__47047\
        );

    \I__10852\ : InMux
    port map (
            O => \N__47097\,
            I => \N__47047\
        );

    \I__10851\ : Span4Mux_v
    port map (
            O => \N__47094\,
            I => \N__47042\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__47089\,
            I => \N__47042\
        );

    \I__10849\ : InMux
    port map (
            O => \N__47088\,
            I => \N__47033\
        );

    \I__10848\ : InMux
    port map (
            O => \N__47087\,
            I => \N__47033\
        );

    \I__10847\ : InMux
    port map (
            O => \N__47086\,
            I => \N__47033\
        );

    \I__10846\ : InMux
    port map (
            O => \N__47085\,
            I => \N__47033\
        );

    \I__10845\ : InMux
    port map (
            O => \N__47084\,
            I => \N__47028\
        );

    \I__10844\ : InMux
    port map (
            O => \N__47083\,
            I => \N__47028\
        );

    \I__10843\ : InMux
    port map (
            O => \N__47080\,
            I => \N__47021\
        );

    \I__10842\ : InMux
    port map (
            O => \N__47079\,
            I => \N__47021\
        );

    \I__10841\ : InMux
    port map (
            O => \N__47078\,
            I => \N__47021\
        );

    \I__10840\ : InMux
    port map (
            O => \N__47077\,
            I => \N__47015\
        );

    \I__10839\ : InMux
    port map (
            O => \N__47076\,
            I => \N__47015\
        );

    \I__10838\ : Span4Mux_v
    port map (
            O => \N__47073\,
            I => \N__47012\
        );

    \I__10837\ : InMux
    port map (
            O => \N__47072\,
            I => \N__46997\
        );

    \I__10836\ : InMux
    port map (
            O => \N__47071\,
            I => \N__46997\
        );

    \I__10835\ : InMux
    port map (
            O => \N__47070\,
            I => \N__46997\
        );

    \I__10834\ : InMux
    port map (
            O => \N__47069\,
            I => \N__46997\
        );

    \I__10833\ : InMux
    port map (
            O => \N__47068\,
            I => \N__46997\
        );

    \I__10832\ : InMux
    port map (
            O => \N__47067\,
            I => \N__46997\
        );

    \I__10831\ : InMux
    port map (
            O => \N__47066\,
            I => \N__46997\
        );

    \I__10830\ : InMux
    port map (
            O => \N__47065\,
            I => \N__46986\
        );

    \I__10829\ : InMux
    port map (
            O => \N__47064\,
            I => \N__46986\
        );

    \I__10828\ : InMux
    port map (
            O => \N__47063\,
            I => \N__46986\
        );

    \I__10827\ : InMux
    port map (
            O => \N__47062\,
            I => \N__46986\
        );

    \I__10826\ : InMux
    port map (
            O => \N__47061\,
            I => \N__46986\
        );

    \I__10825\ : InMux
    port map (
            O => \N__47060\,
            I => \N__46979\
        );

    \I__10824\ : InMux
    port map (
            O => \N__47059\,
            I => \N__46979\
        );

    \I__10823\ : InMux
    port map (
            O => \N__47058\,
            I => \N__46979\
        );

    \I__10822\ : InMux
    port map (
            O => \N__47057\,
            I => \N__46972\
        );

    \I__10821\ : InMux
    port map (
            O => \N__47056\,
            I => \N__46972\
        );

    \I__10820\ : InMux
    port map (
            O => \N__47055\,
            I => \N__46972\
        );

    \I__10819\ : Span4Mux_v
    port map (
            O => \N__47052\,
            I => \N__46959\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__47047\,
            I => \N__46959\
        );

    \I__10817\ : Span4Mux_h
    port map (
            O => \N__47042\,
            I => \N__46959\
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__47033\,
            I => \N__46959\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__47028\,
            I => \N__46959\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__47021\,
            I => \N__46959\
        );

    \I__10813\ : InMux
    port map (
            O => \N__47020\,
            I => \N__46956\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__47015\,
            I => \N__46951\
        );

    \I__10811\ : Span4Mux_h
    port map (
            O => \N__47012\,
            I => \N__46951\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__46997\,
            I => \N__46942\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__46986\,
            I => \N__46942\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__46979\,
            I => \N__46942\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__46972\,
            I => \N__46942\
        );

    \I__10806\ : Span4Mux_v
    port map (
            O => \N__46959\,
            I => \N__46939\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46956\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__10804\ : Odrv4
    port map (
            O => \N__46951\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__10803\ : Odrv12
    port map (
            O => \N__46942\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__10802\ : Odrv4
    port map (
            O => \N__46939\,
            I => \elapsed_time_ns_1_RNI5IV8E1_0_31\
        );

    \I__10801\ : CascadeMux
    port map (
            O => \N__46930\,
            I => \N__46919\
        );

    \I__10800\ : InMux
    port map (
            O => \N__46929\,
            I => \N__46916\
        );

    \I__10799\ : InMux
    port map (
            O => \N__46928\,
            I => \N__46905\
        );

    \I__10798\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46905\
        );

    \I__10797\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46905\
        );

    \I__10796\ : InMux
    port map (
            O => \N__46925\,
            I => \N__46905\
        );

    \I__10795\ : InMux
    port map (
            O => \N__46924\,
            I => \N__46905\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46898\
        );

    \I__10793\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46898\
        );

    \I__10792\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46898\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__46916\,
            I => \phase_controller_inst1.stoper_hc.N_318\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__46905\,
            I => \phase_controller_inst1.stoper_hc.N_318\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__46898\,
            I => \phase_controller_inst1.stoper_hc.N_318\
        );

    \I__10788\ : CascadeMux
    port map (
            O => \N__46891\,
            I => \N__46887\
        );

    \I__10787\ : InMux
    port map (
            O => \N__46890\,
            I => \N__46881\
        );

    \I__10786\ : InMux
    port map (
            O => \N__46887\,
            I => \N__46878\
        );

    \I__10785\ : InMux
    port map (
            O => \N__46886\,
            I => \N__46875\
        );

    \I__10784\ : InMux
    port map (
            O => \N__46885\,
            I => \N__46871\
        );

    \I__10783\ : InMux
    port map (
            O => \N__46884\,
            I => \N__46867\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__46881\,
            I => \N__46864\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46878\,
            I => \N__46861\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__46875\,
            I => \N__46858\
        );

    \I__10779\ : InMux
    port map (
            O => \N__46874\,
            I => \N__46855\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__46871\,
            I => \N__46852\
        );

    \I__10777\ : InMux
    port map (
            O => \N__46870\,
            I => \N__46849\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__46867\,
            I => \N__46838\
        );

    \I__10775\ : Span4Mux_v
    port map (
            O => \N__46864\,
            I => \N__46838\
        );

    \I__10774\ : Span4Mux_v
    port map (
            O => \N__46861\,
            I => \N__46838\
        );

    \I__10773\ : Span4Mux_v
    port map (
            O => \N__46858\,
            I => \N__46838\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__46855\,
            I => \N__46838\
        );

    \I__10771\ : Odrv4
    port map (
            O => \N__46852\,
            I => \elapsed_time_ns_1_RNIDDC6P1_0_14\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46849\,
            I => \elapsed_time_ns_1_RNIDDC6P1_0_14\
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__46838\,
            I => \elapsed_time_ns_1_RNIDDC6P1_0_14\
        );

    \I__10768\ : CascadeMux
    port map (
            O => \N__46831\,
            I => \N__46819\
        );

    \I__10767\ : CascadeMux
    port map (
            O => \N__46830\,
            I => \N__46816\
        );

    \I__10766\ : CascadeMux
    port map (
            O => \N__46829\,
            I => \N__46813\
        );

    \I__10765\ : InMux
    port map (
            O => \N__46828\,
            I => \N__46807\
        );

    \I__10764\ : CascadeMux
    port map (
            O => \N__46827\,
            I => \N__46796\
        );

    \I__10763\ : InMux
    port map (
            O => \N__46826\,
            I => \N__46791\
        );

    \I__10762\ : InMux
    port map (
            O => \N__46825\,
            I => \N__46776\
        );

    \I__10761\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46776\
        );

    \I__10760\ : InMux
    port map (
            O => \N__46823\,
            I => \N__46776\
        );

    \I__10759\ : InMux
    port map (
            O => \N__46822\,
            I => \N__46776\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46819\,
            I => \N__46776\
        );

    \I__10757\ : InMux
    port map (
            O => \N__46816\,
            I => \N__46776\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46776\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46812\,
            I => \N__46773\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46811\,
            I => \N__46768\
        );

    \I__10753\ : InMux
    port map (
            O => \N__46810\,
            I => \N__46768\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__46807\,
            I => \N__46765\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46806\,
            I => \N__46754\
        );

    \I__10750\ : InMux
    port map (
            O => \N__46805\,
            I => \N__46754\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46804\,
            I => \N__46754\
        );

    \I__10748\ : InMux
    port map (
            O => \N__46803\,
            I => \N__46754\
        );

    \I__10747\ : InMux
    port map (
            O => \N__46802\,
            I => \N__46754\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46801\,
            I => \N__46751\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46800\,
            I => \N__46748\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46799\,
            I => \N__46742\
        );

    \I__10743\ : InMux
    port map (
            O => \N__46796\,
            I => \N__46735\
        );

    \I__10742\ : InMux
    port map (
            O => \N__46795\,
            I => \N__46735\
        );

    \I__10741\ : InMux
    port map (
            O => \N__46794\,
            I => \N__46735\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__46791\,
            I => \N__46732\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__46776\,
            I => \N__46729\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__46773\,
            I => \N__46726\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__46768\,
            I => \N__46719\
        );

    \I__10736\ : Span4Mux_v
    port map (
            O => \N__46765\,
            I => \N__46719\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__46754\,
            I => \N__46719\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__46751\,
            I => \N__46714\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__46748\,
            I => \N__46714\
        );

    \I__10732\ : InMux
    port map (
            O => \N__46747\,
            I => \N__46709\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46746\,
            I => \N__46709\
        );

    \I__10730\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46706\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__46742\,
            I => \N__46699\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__46735\,
            I => \N__46699\
        );

    \I__10727\ : Span4Mux_h
    port map (
            O => \N__46732\,
            I => \N__46699\
        );

    \I__10726\ : Span4Mux_v
    port map (
            O => \N__46729\,
            I => \N__46694\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__46726\,
            I => \N__46694\
        );

    \I__10724\ : Span4Mux_v
    port map (
            O => \N__46719\,
            I => \N__46687\
        );

    \I__10723\ : Span4Mux_v
    port map (
            O => \N__46714\,
            I => \N__46687\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__46709\,
            I => \N__46687\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__46706\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__10720\ : Odrv4
    port map (
            O => \N__46699\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__10719\ : Odrv4
    port map (
            O => \N__46694\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__10718\ : Odrv4
    port map (
            O => \N__46687\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\
        );

    \I__10717\ : CascadeMux
    port map (
            O => \N__46678\,
            I => \N__46675\
        );

    \I__10716\ : InMux
    port map (
            O => \N__46675\,
            I => \N__46672\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__46672\,
            I => \N__46669\
        );

    \I__10714\ : Odrv12
    port map (
            O => \N__46669\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__10713\ : InMux
    port map (
            O => \N__46666\,
            I => \N__46660\
        );

    \I__10712\ : InMux
    port map (
            O => \N__46665\,
            I => \N__46657\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46664\,
            I => \N__46653\
        );

    \I__10710\ : InMux
    port map (
            O => \N__46663\,
            I => \N__46650\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__46660\,
            I => \N__46647\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__46657\,
            I => \N__46644\
        );

    \I__10707\ : CascadeMux
    port map (
            O => \N__46656\,
            I => \N__46640\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__46653\,
            I => \N__46635\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__46650\,
            I => \N__46635\
        );

    \I__10704\ : Span4Mux_v
    port map (
            O => \N__46647\,
            I => \N__46632\
        );

    \I__10703\ : Sp12to4
    port map (
            O => \N__46644\,
            I => \N__46629\
        );

    \I__10702\ : InMux
    port map (
            O => \N__46643\,
            I => \N__46626\
        );

    \I__10701\ : InMux
    port map (
            O => \N__46640\,
            I => \N__46623\
        );

    \I__10700\ : Span4Mux_v
    port map (
            O => \N__46635\,
            I => \N__46618\
        );

    \I__10699\ : Span4Mux_h
    port map (
            O => \N__46632\,
            I => \N__46618\
        );

    \I__10698\ : Span12Mux_h
    port map (
            O => \N__46629\,
            I => \N__46615\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__46626\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__46623\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__10695\ : Odrv4
    port map (
            O => \N__46618\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__10694\ : Odrv12
    port map (
            O => \N__46615\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__10693\ : CascadeMux
    port map (
            O => \N__46606\,
            I => \N__46603\
        );

    \I__10692\ : InMux
    port map (
            O => \N__46603\,
            I => \N__46600\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__46600\,
            I => \N__46595\
        );

    \I__10690\ : InMux
    port map (
            O => \N__46599\,
            I => \N__46592\
        );

    \I__10689\ : InMux
    port map (
            O => \N__46598\,
            I => \N__46589\
        );

    \I__10688\ : Span4Mux_h
    port map (
            O => \N__46595\,
            I => \N__46584\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__46592\,
            I => \N__46581\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__46589\,
            I => \N__46578\
        );

    \I__10685\ : InMux
    port map (
            O => \N__46588\,
            I => \N__46575\
        );

    \I__10684\ : InMux
    port map (
            O => \N__46587\,
            I => \N__46572\
        );

    \I__10683\ : Span4Mux_v
    port map (
            O => \N__46584\,
            I => \N__46569\
        );

    \I__10682\ : Span4Mux_h
    port map (
            O => \N__46581\,
            I => \N__46564\
        );

    \I__10681\ : Span4Mux_h
    port map (
            O => \N__46578\,
            I => \N__46564\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__46575\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__46572\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__10678\ : Odrv4
    port map (
            O => \N__46569\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__10677\ : Odrv4
    port map (
            O => \N__46564\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__10676\ : IoInMux
    port map (
            O => \N__46555\,
            I => \N__46552\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__46552\,
            I => \N__46549\
        );

    \I__10674\ : Span4Mux_s1_v
    port map (
            O => \N__46549\,
            I => \N__46546\
        );

    \I__10673\ : Span4Mux_v
    port map (
            O => \N__46546\,
            I => \N__46542\
        );

    \I__10672\ : InMux
    port map (
            O => \N__46545\,
            I => \N__46539\
        );

    \I__10671\ : Odrv4
    port map (
            O => \N__46542\,
            I => \T12_c\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__46539\,
            I => \T12_c\
        );

    \I__10669\ : CascadeMux
    port map (
            O => \N__46534\,
            I => \N__46530\
        );

    \I__10668\ : InMux
    port map (
            O => \N__46533\,
            I => \N__46527\
        );

    \I__10667\ : InMux
    port map (
            O => \N__46530\,
            I => \N__46524\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__46527\,
            I => \N__46521\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__46524\,
            I => \N__46517\
        );

    \I__10664\ : Span4Mux_v
    port map (
            O => \N__46521\,
            I => \N__46514\
        );

    \I__10663\ : InMux
    port map (
            O => \N__46520\,
            I => \N__46511\
        );

    \I__10662\ : Span4Mux_v
    port map (
            O => \N__46517\,
            I => \N__46508\
        );

    \I__10661\ : Odrv4
    port map (
            O => \N__46514\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__46511\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10659\ : Odrv4
    port map (
            O => \N__46508\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10658\ : CascadeMux
    port map (
            O => \N__46501\,
            I => \N__46498\
        );

    \I__10657\ : InMux
    port map (
            O => \N__46498\,
            I => \N__46495\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__46495\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__10655\ : InMux
    port map (
            O => \N__46492\,
            I => \N__46489\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__46489\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__10653\ : InMux
    port map (
            O => \N__46486\,
            I => \N__46483\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__46483\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__10651\ : CascadeMux
    port map (
            O => \N__46480\,
            I => \N__46477\
        );

    \I__10650\ : InMux
    port map (
            O => \N__46477\,
            I => \N__46474\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__46474\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__10648\ : InMux
    port map (
            O => \N__46471\,
            I => \N__46468\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__46468\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__10646\ : InMux
    port map (
            O => \N__46465\,
            I => \N__46462\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__46462\,
            I => \N__46459\
        );

    \I__10644\ : Odrv4
    port map (
            O => \N__46459\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__10643\ : CascadeMux
    port map (
            O => \N__46456\,
            I => \N__46453\
        );

    \I__10642\ : InMux
    port map (
            O => \N__46453\,
            I => \N__46450\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__46450\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__10640\ : InMux
    port map (
            O => \N__46447\,
            I => \N__46444\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__46444\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__10638\ : CascadeMux
    port map (
            O => \N__46441\,
            I => \N__46438\
        );

    \I__10637\ : InMux
    port map (
            O => \N__46438\,
            I => \N__46435\
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__46435\,
            I => \N__46432\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__46432\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__10634\ : InMux
    port map (
            O => \N__46429\,
            I => \N__46426\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__46426\,
            I => \N__46423\
        );

    \I__10632\ : Odrv4
    port map (
            O => \N__46423\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__46420\,
            I => \N__46417\
        );

    \I__10630\ : InMux
    port map (
            O => \N__46417\,
            I => \N__46414\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__46414\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__10628\ : InMux
    port map (
            O => \N__46411\,
            I => \N__46408\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__46408\,
            I => \N__46405\
        );

    \I__10626\ : Odrv12
    port map (
            O => \N__46405\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__10625\ : CascadeMux
    port map (
            O => \N__46402\,
            I => \N__46399\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46399\,
            I => \N__46396\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__46396\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__10622\ : InMux
    port map (
            O => \N__46393\,
            I => \N__46390\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__46390\,
            I => \N__46387\
        );

    \I__10620\ : Span4Mux_v
    port map (
            O => \N__46387\,
            I => \N__46384\
        );

    \I__10619\ : Odrv4
    port map (
            O => \N__46384\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__10618\ : CascadeMux
    port map (
            O => \N__46381\,
            I => \N__46378\
        );

    \I__10617\ : InMux
    port map (
            O => \N__46378\,
            I => \N__46375\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__46375\,
            I => \N__46372\
        );

    \I__10615\ : Odrv4
    port map (
            O => \N__46372\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__10614\ : InMux
    port map (
            O => \N__46369\,
            I => \N__46366\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__46366\,
            I => \N__46363\
        );

    \I__10612\ : Span4Mux_v
    port map (
            O => \N__46363\,
            I => \N__46360\
        );

    \I__10611\ : Span4Mux_h
    port map (
            O => \N__46360\,
            I => \N__46357\
        );

    \I__10610\ : Odrv4
    port map (
            O => \N__46357\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__10609\ : CascadeMux
    port map (
            O => \N__46354\,
            I => \N__46351\
        );

    \I__10608\ : InMux
    port map (
            O => \N__46351\,
            I => \N__46348\
        );

    \I__10607\ : LocalMux
    port map (
            O => \N__46348\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__10606\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46342\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__46342\,
            I => \N__46339\
        );

    \I__10604\ : Span4Mux_v
    port map (
            O => \N__46339\,
            I => \N__46336\
        );

    \I__10603\ : Span4Mux_h
    port map (
            O => \N__46336\,
            I => \N__46333\
        );

    \I__10602\ : Odrv4
    port map (
            O => \N__46333\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__10601\ : CascadeMux
    port map (
            O => \N__46330\,
            I => \N__46327\
        );

    \I__10600\ : InMux
    port map (
            O => \N__46327\,
            I => \N__46324\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__46324\,
            I => \N__46321\
        );

    \I__10598\ : Odrv4
    port map (
            O => \N__46321\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__10597\ : InMux
    port map (
            O => \N__46318\,
            I => \N__46315\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__46315\,
            I => \N__46312\
        );

    \I__10595\ : Odrv12
    port map (
            O => \N__46312\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__10594\ : CascadeMux
    port map (
            O => \N__46309\,
            I => \N__46306\
        );

    \I__10593\ : InMux
    port map (
            O => \N__46306\,
            I => \N__46303\
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__46303\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__10591\ : InMux
    port map (
            O => \N__46300\,
            I => \N__46297\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__46297\,
            I => \N__46294\
        );

    \I__10589\ : Odrv4
    port map (
            O => \N__46294\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__10588\ : CascadeMux
    port map (
            O => \N__46291\,
            I => \N__46288\
        );

    \I__10587\ : InMux
    port map (
            O => \N__46288\,
            I => \N__46285\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__46285\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__10585\ : InMux
    port map (
            O => \N__46282\,
            I => \N__46279\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__46279\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__10583\ : CascadeMux
    port map (
            O => \N__46276\,
            I => \N__46273\
        );

    \I__10582\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46270\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__46270\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__10580\ : InMux
    port map (
            O => \N__46267\,
            I => \N__46264\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__46264\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__10578\ : CascadeMux
    port map (
            O => \N__46261\,
            I => \N__46258\
        );

    \I__10577\ : InMux
    port map (
            O => \N__46258\,
            I => \N__46255\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__46255\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__10575\ : CascadeMux
    port map (
            O => \N__46252\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__10574\ : CascadeMux
    port map (
            O => \N__46249\,
            I => \N__46246\
        );

    \I__10573\ : InMux
    port map (
            O => \N__46246\,
            I => \N__46240\
        );

    \I__10572\ : InMux
    port map (
            O => \N__46245\,
            I => \N__46240\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__46240\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__10570\ : CascadeMux
    port map (
            O => \N__46237\,
            I => \N__46234\
        );

    \I__10569\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46228\
        );

    \I__10568\ : InMux
    port map (
            O => \N__46233\,
            I => \N__46228\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__46228\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__10566\ : CascadeMux
    port map (
            O => \N__46225\,
            I => \N__46222\
        );

    \I__10565\ : InMux
    port map (
            O => \N__46222\,
            I => \N__46215\
        );

    \I__10564\ : InMux
    port map (
            O => \N__46221\,
            I => \N__46206\
        );

    \I__10563\ : InMux
    port map (
            O => \N__46220\,
            I => \N__46206\
        );

    \I__10562\ : InMux
    port map (
            O => \N__46219\,
            I => \N__46206\
        );

    \I__10561\ : InMux
    port map (
            O => \N__46218\,
            I => \N__46206\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__46215\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__46206\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__10558\ : CascadeMux
    port map (
            O => \N__46201\,
            I => \N__46198\
        );

    \I__10557\ : InMux
    port map (
            O => \N__46198\,
            I => \N__46194\
        );

    \I__10556\ : CascadeMux
    port map (
            O => \N__46197\,
            I => \N__46191\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46194\,
            I => \N__46187\
        );

    \I__10554\ : InMux
    port map (
            O => \N__46191\,
            I => \N__46182\
        );

    \I__10553\ : InMux
    port map (
            O => \N__46190\,
            I => \N__46182\
        );

    \I__10552\ : Span4Mux_v
    port map (
            O => \N__46187\,
            I => \N__46178\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__46182\,
            I => \N__46175\
        );

    \I__10550\ : InMux
    port map (
            O => \N__46181\,
            I => \N__46172\
        );

    \I__10549\ : Span4Mux_h
    port map (
            O => \N__46178\,
            I => \N__46169\
        );

    \I__10548\ : Span4Mux_v
    port map (
            O => \N__46175\,
            I => \N__46166\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__46172\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__10546\ : Odrv4
    port map (
            O => \N__46169\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__10545\ : Odrv4
    port map (
            O => \N__46166\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__10544\ : InMux
    port map (
            O => \N__46159\,
            I => \N__46153\
        );

    \I__10543\ : InMux
    port map (
            O => \N__46158\,
            I => \N__46153\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__46153\,
            I => \N__46148\
        );

    \I__10541\ : InMux
    port map (
            O => \N__46152\,
            I => \N__46143\
        );

    \I__10540\ : InMux
    port map (
            O => \N__46151\,
            I => \N__46143\
        );

    \I__10539\ : Span4Mux_v
    port map (
            O => \N__46148\,
            I => \N__46140\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__46143\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__10537\ : Odrv4
    port map (
            O => \N__46140\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__10536\ : InMux
    port map (
            O => \N__46135\,
            I => \N__46132\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__46132\,
            I => \N__46129\
        );

    \I__10534\ : Span4Mux_v
    port map (
            O => \N__46129\,
            I => \N__46122\
        );

    \I__10533\ : InMux
    port map (
            O => \N__46128\,
            I => \N__46113\
        );

    \I__10532\ : InMux
    port map (
            O => \N__46127\,
            I => \N__46113\
        );

    \I__10531\ : InMux
    port map (
            O => \N__46126\,
            I => \N__46113\
        );

    \I__10530\ : InMux
    port map (
            O => \N__46125\,
            I => \N__46113\
        );

    \I__10529\ : Odrv4
    port map (
            O => \N__46122\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__46113\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__10527\ : InMux
    port map (
            O => \N__46108\,
            I => \N__46105\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__46105\,
            I => \N__46102\
        );

    \I__10525\ : Odrv12
    port map (
            O => \N__46102\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__10524\ : CascadeMux
    port map (
            O => \N__46099\,
            I => \N__46096\
        );

    \I__10523\ : InMux
    port map (
            O => \N__46096\,
            I => \N__46093\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__46093\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__10521\ : InMux
    port map (
            O => \N__46090\,
            I => \N__46087\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__46087\,
            I => \N__46084\
        );

    \I__10519\ : Span4Mux_h
    port map (
            O => \N__46084\,
            I => \N__46081\
        );

    \I__10518\ : Odrv4
    port map (
            O => \N__46081\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__10517\ : CascadeMux
    port map (
            O => \N__46078\,
            I => \N__46075\
        );

    \I__10516\ : InMux
    port map (
            O => \N__46075\,
            I => \N__46072\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__46072\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__10514\ : InMux
    port map (
            O => \N__46069\,
            I => \N__46066\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__46066\,
            I => \N__46063\
        );

    \I__10512\ : Span4Mux_h
    port map (
            O => \N__46063\,
            I => \N__46060\
        );

    \I__10511\ : Odrv4
    port map (
            O => \N__46060\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__10510\ : CascadeMux
    port map (
            O => \N__46057\,
            I => \N__46054\
        );

    \I__10509\ : InMux
    port map (
            O => \N__46054\,
            I => \N__46051\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__46051\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__10507\ : InMux
    port map (
            O => \N__46048\,
            I => \N__46044\
        );

    \I__10506\ : InMux
    port map (
            O => \N__46047\,
            I => \N__46041\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__46044\,
            I => \N__46038\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__46041\,
            I => \N__46035\
        );

    \I__10503\ : Span4Mux_h
    port map (
            O => \N__46038\,
            I => \N__46032\
        );

    \I__10502\ : Odrv4
    port map (
            O => \N__46035\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__10501\ : Odrv4
    port map (
            O => \N__46032\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__10500\ : CascadeMux
    port map (
            O => \N__46027\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_\
        );

    \I__10499\ : InMux
    port map (
            O => \N__46024\,
            I => \N__46020\
        );

    \I__10498\ : InMux
    port map (
            O => \N__46023\,
            I => \N__46017\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__46020\,
            I => \N__46008\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__46017\,
            I => \N__46008\
        );

    \I__10495\ : InMux
    port map (
            O => \N__46016\,
            I => \N__46005\
        );

    \I__10494\ : InMux
    port map (
            O => \N__46015\,
            I => \N__46001\
        );

    \I__10493\ : InMux
    port map (
            O => \N__46014\,
            I => \N__45997\
        );

    \I__10492\ : InMux
    port map (
            O => \N__46013\,
            I => \N__45994\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__46008\,
            I => \N__45991\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__46005\,
            I => \N__45988\
        );

    \I__10489\ : InMux
    port map (
            O => \N__46004\,
            I => \N__45985\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__46001\,
            I => \N__45982\
        );

    \I__10487\ : InMux
    port map (
            O => \N__46000\,
            I => \N__45979\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__45997\,
            I => \delay_measurement_inst.delay_hc_timer.N_344_i\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45994\,
            I => \delay_measurement_inst.delay_hc_timer.N_344_i\
        );

    \I__10484\ : Odrv4
    port map (
            O => \N__45991\,
            I => \delay_measurement_inst.delay_hc_timer.N_344_i\
        );

    \I__10483\ : Odrv4
    port map (
            O => \N__45988\,
            I => \delay_measurement_inst.delay_hc_timer.N_344_i\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__45985\,
            I => \delay_measurement_inst.delay_hc_timer.N_344_i\
        );

    \I__10481\ : Odrv12
    port map (
            O => \N__45982\,
            I => \delay_measurement_inst.delay_hc_timer.N_344_i\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__45979\,
            I => \delay_measurement_inst.delay_hc_timer.N_344_i\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45964\,
            I => \N__45961\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__45961\,
            I => \N__45955\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45960\,
            I => \N__45950\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45959\,
            I => \N__45950\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45958\,
            I => \N__45947\
        );

    \I__10474\ : Span12Mux_v
    port map (
            O => \N__45955\,
            I => \N__45942\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__45950\,
            I => \N__45942\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__45947\,
            I => \elapsed_time_ns_1_RNIUE3CP1_0_6\
        );

    \I__10471\ : Odrv12
    port map (
            O => \N__45942\,
            I => \elapsed_time_ns_1_RNIUE3CP1_0_6\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45937\,
            I => \N__45933\
        );

    \I__10469\ : CascadeMux
    port map (
            O => \N__45936\,
            I => \N__45930\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__45933\,
            I => \N__45923\
        );

    \I__10467\ : InMux
    port map (
            O => \N__45930\,
            I => \N__45919\
        );

    \I__10466\ : InMux
    port map (
            O => \N__45929\,
            I => \N__45916\
        );

    \I__10465\ : CascadeMux
    port map (
            O => \N__45928\,
            I => \N__45912\
        );

    \I__10464\ : CascadeMux
    port map (
            O => \N__45927\,
            I => \N__45908\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45926\,
            I => \N__45899\
        );

    \I__10462\ : Span4Mux_v
    port map (
            O => \N__45923\,
            I => \N__45896\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45922\,
            I => \N__45893\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__45919\,
            I => \N__45888\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__45916\,
            I => \N__45888\
        );

    \I__10458\ : InMux
    port map (
            O => \N__45915\,
            I => \N__45881\
        );

    \I__10457\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45881\
        );

    \I__10456\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45881\
        );

    \I__10455\ : InMux
    port map (
            O => \N__45908\,
            I => \N__45878\
        );

    \I__10454\ : CascadeMux
    port map (
            O => \N__45907\,
            I => \N__45875\
        );

    \I__10453\ : CascadeMux
    port map (
            O => \N__45906\,
            I => \N__45869\
        );

    \I__10452\ : CascadeMux
    port map (
            O => \N__45905\,
            I => \N__45865\
        );

    \I__10451\ : CascadeMux
    port map (
            O => \N__45904\,
            I => \N__45862\
        );

    \I__10450\ : InMux
    port map (
            O => \N__45903\,
            I => \N__45855\
        );

    \I__10449\ : InMux
    port map (
            O => \N__45902\,
            I => \N__45855\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__45899\,
            I => \N__45848\
        );

    \I__10447\ : Span4Mux_h
    port map (
            O => \N__45896\,
            I => \N__45848\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45893\,
            I => \N__45848\
        );

    \I__10445\ : Span4Mux_h
    port map (
            O => \N__45888\,
            I => \N__45841\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__45881\,
            I => \N__45841\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__45878\,
            I => \N__45841\
        );

    \I__10442\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45830\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45830\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45830\
        );

    \I__10439\ : InMux
    port map (
            O => \N__45872\,
            I => \N__45830\
        );

    \I__10438\ : InMux
    port map (
            O => \N__45869\,
            I => \N__45830\
        );

    \I__10437\ : InMux
    port map (
            O => \N__45868\,
            I => \N__45819\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45865\,
            I => \N__45819\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45862\,
            I => \N__45819\
        );

    \I__10434\ : InMux
    port map (
            O => \N__45861\,
            I => \N__45819\
        );

    \I__10433\ : InMux
    port map (
            O => \N__45860\,
            I => \N__45819\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__45855\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__10431\ : Odrv4
    port map (
            O => \N__45848\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__10430\ : Odrv4
    port map (
            O => \N__45841\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__45830\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45819\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\
        );

    \I__10427\ : InMux
    port map (
            O => \N__45808\,
            I => \N__45805\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__45805\,
            I => \N__45802\
        );

    \I__10425\ : Span4Mux_h
    port map (
            O => \N__45802\,
            I => \N__45798\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45801\,
            I => \N__45795\
        );

    \I__10423\ : Odrv4
    port map (
            O => \N__45798\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__45795\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10421\ : CascadeMux
    port map (
            O => \N__45790\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15_cascade_\
        );

    \I__10420\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45783\
        );

    \I__10419\ : InMux
    port map (
            O => \N__45786\,
            I => \N__45780\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__45783\,
            I => \N__45774\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__45780\,
            I => \N__45774\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45779\,
            I => \N__45771\
        );

    \I__10415\ : Span4Mux_v
    port map (
            O => \N__45774\,
            I => \N__45768\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__45771\,
            I => \N__45765\
        );

    \I__10413\ : Span4Mux_h
    port map (
            O => \N__45768\,
            I => \N__45762\
        );

    \I__10412\ : Odrv4
    port map (
            O => \N__45765\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\
        );

    \I__10411\ : Odrv4
    port map (
            O => \N__45762\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\
        );

    \I__10410\ : InMux
    port map (
            O => \N__45757\,
            I => \N__45753\
        );

    \I__10409\ : InMux
    port map (
            O => \N__45756\,
            I => \N__45750\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__45753\,
            I => \N__45747\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__45750\,
            I => \N__45744\
        );

    \I__10406\ : Span4Mux_h
    port map (
            O => \N__45747\,
            I => \N__45739\
        );

    \I__10405\ : Span4Mux_v
    port map (
            O => \N__45744\,
            I => \N__45739\
        );

    \I__10404\ : Odrv4
    port map (
            O => \N__45739\,
            I => \phase_controller_inst1.stoper_hc.N_269_iZ0Z_1\
        );

    \I__10403\ : CascadeMux
    port map (
            O => \N__45736\,
            I => \N__45732\
        );

    \I__10402\ : InMux
    port map (
            O => \N__45735\,
            I => \N__45727\
        );

    \I__10401\ : InMux
    port map (
            O => \N__45732\,
            I => \N__45724\
        );

    \I__10400\ : InMux
    port map (
            O => \N__45731\,
            I => \N__45721\
        );

    \I__10399\ : CascadeMux
    port map (
            O => \N__45730\,
            I => \N__45718\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__45727\,
            I => \N__45714\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__45724\,
            I => \N__45709\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__45721\,
            I => \N__45709\
        );

    \I__10395\ : InMux
    port map (
            O => \N__45718\,
            I => \N__45706\
        );

    \I__10394\ : CascadeMux
    port map (
            O => \N__45717\,
            I => \N__45702\
        );

    \I__10393\ : Span4Mux_v
    port map (
            O => \N__45714\,
            I => \N__45694\
        );

    \I__10392\ : Span4Mux_v
    port map (
            O => \N__45709\,
            I => \N__45694\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__45706\,
            I => \N__45694\
        );

    \I__10390\ : InMux
    port map (
            O => \N__45705\,
            I => \N__45691\
        );

    \I__10389\ : InMux
    port map (
            O => \N__45702\,
            I => \N__45686\
        );

    \I__10388\ : InMux
    port map (
            O => \N__45701\,
            I => \N__45686\
        );

    \I__10387\ : Span4Mux_h
    port map (
            O => \N__45694\,
            I => \N__45683\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__45691\,
            I => \N__45680\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__45686\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15\
        );

    \I__10384\ : Odrv4
    port map (
            O => \N__45683\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15\
        );

    \I__10383\ : Odrv12
    port map (
            O => \N__45680\,
            I => \elapsed_time_ns_1_RNI7IT8E1_0_15\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45673\,
            I => \N__45669\
        );

    \I__10381\ : InMux
    port map (
            O => \N__45672\,
            I => \N__45665\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__45669\,
            I => \N__45662\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45659\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__45665\,
            I => \N__45656\
        );

    \I__10377\ : Span4Mux_v
    port map (
            O => \N__45662\,
            I => \N__45649\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__45659\,
            I => \N__45649\
        );

    \I__10375\ : Span4Mux_h
    port map (
            O => \N__45656\,
            I => \N__45646\
        );

    \I__10374\ : InMux
    port map (
            O => \N__45655\,
            I => \N__45641\
        );

    \I__10373\ : InMux
    port map (
            O => \N__45654\,
            I => \N__45641\
        );

    \I__10372\ : Span4Mux_h
    port map (
            O => \N__45649\,
            I => \N__45638\
        );

    \I__10371\ : Odrv4
    port map (
            O => \N__45646\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__45641\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__10369\ : Odrv4
    port map (
            O => \N__45638\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\
        );

    \I__10368\ : CascadeMux
    port map (
            O => \N__45631\,
            I => \N__45627\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45624\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45627\,
            I => \N__45621\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__45624\,
            I => \N__45618\
        );

    \I__10364\ : LocalMux
    port map (
            O => \N__45621\,
            I => \N__45615\
        );

    \I__10363\ : Odrv4
    port map (
            O => \N__45618\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__10362\ : Odrv12
    port map (
            O => \N__45615\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__10361\ : CascadeMux
    port map (
            O => \N__45610\,
            I => \N__45606\
        );

    \I__10360\ : InMux
    port map (
            O => \N__45609\,
            I => \N__45603\
        );

    \I__10359\ : InMux
    port map (
            O => \N__45606\,
            I => \N__45599\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__45603\,
            I => \N__45596\
        );

    \I__10357\ : CascadeMux
    port map (
            O => \N__45602\,
            I => \N__45593\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__45599\,
            I => \N__45590\
        );

    \I__10355\ : Span4Mux_v
    port map (
            O => \N__45596\,
            I => \N__45585\
        );

    \I__10354\ : InMux
    port map (
            O => \N__45593\,
            I => \N__45582\
        );

    \I__10353\ : Span4Mux_h
    port map (
            O => \N__45590\,
            I => \N__45579\
        );

    \I__10352\ : InMux
    port map (
            O => \N__45589\,
            I => \N__45576\
        );

    \I__10351\ : InMux
    port map (
            O => \N__45588\,
            I => \N__45573\
        );

    \I__10350\ : Odrv4
    port map (
            O => \N__45585\,
            I => \elapsed_time_ns_1_RNI1I3CP1_0_9\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__45582\,
            I => \elapsed_time_ns_1_RNI1I3CP1_0_9\
        );

    \I__10348\ : Odrv4
    port map (
            O => \N__45579\,
            I => \elapsed_time_ns_1_RNI1I3CP1_0_9\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__45576\,
            I => \elapsed_time_ns_1_RNI1I3CP1_0_9\
        );

    \I__10346\ : LocalMux
    port map (
            O => \N__45573\,
            I => \elapsed_time_ns_1_RNI1I3CP1_0_9\
        );

    \I__10345\ : CascadeMux
    port map (
            O => \N__45562\,
            I => \N__45557\
        );

    \I__10344\ : InMux
    port map (
            O => \N__45561\,
            I => \N__45553\
        );

    \I__10343\ : InMux
    port map (
            O => \N__45560\,
            I => \N__45540\
        );

    \I__10342\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45540\
        );

    \I__10341\ : CascadeMux
    port map (
            O => \N__45556\,
            I => \N__45537\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__45553\,
            I => \N__45534\
        );

    \I__10339\ : CascadeMux
    port map (
            O => \N__45552\,
            I => \N__45531\
        );

    \I__10338\ : CascadeMux
    port map (
            O => \N__45551\,
            I => \N__45528\
        );

    \I__10337\ : CascadeMux
    port map (
            O => \N__45550\,
            I => \N__45525\
        );

    \I__10336\ : CascadeMux
    port map (
            O => \N__45549\,
            I => \N__45521\
        );

    \I__10335\ : InMux
    port map (
            O => \N__45548\,
            I => \N__45518\
        );

    \I__10334\ : InMux
    port map (
            O => \N__45547\,
            I => \N__45515\
        );

    \I__10333\ : InMux
    port map (
            O => \N__45546\,
            I => \N__45508\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45545\,
            I => \N__45505\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__45540\,
            I => \N__45502\
        );

    \I__10330\ : InMux
    port map (
            O => \N__45537\,
            I => \N__45499\
        );

    \I__10329\ : Span4Mux_v
    port map (
            O => \N__45534\,
            I => \N__45496\
        );

    \I__10328\ : InMux
    port map (
            O => \N__45531\,
            I => \N__45491\
        );

    \I__10327\ : InMux
    port map (
            O => \N__45528\,
            I => \N__45491\
        );

    \I__10326\ : InMux
    port map (
            O => \N__45525\,
            I => \N__45486\
        );

    \I__10325\ : InMux
    port map (
            O => \N__45524\,
            I => \N__45486\
        );

    \I__10324\ : InMux
    port map (
            O => \N__45521\,
            I => \N__45483\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__45518\,
            I => \N__45478\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__45515\,
            I => \N__45478\
        );

    \I__10321\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45471\
        );

    \I__10320\ : InMux
    port map (
            O => \N__45513\,
            I => \N__45471\
        );

    \I__10319\ : InMux
    port map (
            O => \N__45512\,
            I => \N__45471\
        );

    \I__10318\ : CascadeMux
    port map (
            O => \N__45511\,
            I => \N__45467\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__45508\,
            I => \N__45450\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__45505\,
            I => \N__45450\
        );

    \I__10315\ : Span4Mux_h
    port map (
            O => \N__45502\,
            I => \N__45447\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__45499\,
            I => \N__45436\
        );

    \I__10313\ : Span4Mux_h
    port map (
            O => \N__45496\,
            I => \N__45436\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__45491\,
            I => \N__45436\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__45486\,
            I => \N__45436\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__45483\,
            I => \N__45436\
        );

    \I__10309\ : Span4Mux_h
    port map (
            O => \N__45478\,
            I => \N__45431\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__45471\,
            I => \N__45431\
        );

    \I__10307\ : InMux
    port map (
            O => \N__45470\,
            I => \N__45428\
        );

    \I__10306\ : InMux
    port map (
            O => \N__45467\,
            I => \N__45425\
        );

    \I__10305\ : InMux
    port map (
            O => \N__45466\,
            I => \N__45420\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45465\,
            I => \N__45420\
        );

    \I__10303\ : InMux
    port map (
            O => \N__45464\,
            I => \N__45409\
        );

    \I__10302\ : InMux
    port map (
            O => \N__45463\,
            I => \N__45409\
        );

    \I__10301\ : InMux
    port map (
            O => \N__45462\,
            I => \N__45409\
        );

    \I__10300\ : InMux
    port map (
            O => \N__45461\,
            I => \N__45409\
        );

    \I__10299\ : InMux
    port map (
            O => \N__45460\,
            I => \N__45409\
        );

    \I__10298\ : InMux
    port map (
            O => \N__45459\,
            I => \N__45398\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45398\
        );

    \I__10296\ : InMux
    port map (
            O => \N__45457\,
            I => \N__45398\
        );

    \I__10295\ : InMux
    port map (
            O => \N__45456\,
            I => \N__45398\
        );

    \I__10294\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45398\
        );

    \I__10293\ : Odrv12
    port map (
            O => \N__45450\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk\
        );

    \I__10292\ : Odrv4
    port map (
            O => \N__45447\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk\
        );

    \I__10291\ : Odrv4
    port map (
            O => \N__45436\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk\
        );

    \I__10290\ : Odrv4
    port map (
            O => \N__45431\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__45428\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__45425\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__45420\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__45409\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__45398\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk\
        );

    \I__10284\ : CascadeMux
    port map (
            O => \N__45379\,
            I => \N__45376\
        );

    \I__10283\ : InMux
    port map (
            O => \N__45376\,
            I => \N__45371\
        );

    \I__10282\ : InMux
    port map (
            O => \N__45375\,
            I => \N__45365\
        );

    \I__10281\ : InMux
    port map (
            O => \N__45374\,
            I => \N__45365\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__45371\,
            I => \N__45361\
        );

    \I__10279\ : InMux
    port map (
            O => \N__45370\,
            I => \N__45358\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45365\,
            I => \N__45355\
        );

    \I__10277\ : CascadeMux
    port map (
            O => \N__45364\,
            I => \N__45349\
        );

    \I__10276\ : Span4Mux_h
    port map (
            O => \N__45361\,
            I => \N__45343\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__45358\,
            I => \N__45343\
        );

    \I__10274\ : Span4Mux_h
    port map (
            O => \N__45355\,
            I => \N__45340\
        );

    \I__10273\ : InMux
    port map (
            O => \N__45354\,
            I => \N__45337\
        );

    \I__10272\ : CascadeMux
    port map (
            O => \N__45353\,
            I => \N__45329\
        );

    \I__10271\ : CascadeMux
    port map (
            O => \N__45352\,
            I => \N__45326\
        );

    \I__10270\ : InMux
    port map (
            O => \N__45349\,
            I => \N__45323\
        );

    \I__10269\ : InMux
    port map (
            O => \N__45348\,
            I => \N__45320\
        );

    \I__10268\ : Span4Mux_v
    port map (
            O => \N__45343\,
            I => \N__45317\
        );

    \I__10267\ : Span4Mux_v
    port map (
            O => \N__45340\,
            I => \N__45306\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__45337\,
            I => \N__45306\
        );

    \I__10265\ : CascadeMux
    port map (
            O => \N__45336\,
            I => \N__45303\
        );

    \I__10264\ : CascadeMux
    port map (
            O => \N__45335\,
            I => \N__45300\
        );

    \I__10263\ : CascadeMux
    port map (
            O => \N__45334\,
            I => \N__45297\
        );

    \I__10262\ : InMux
    port map (
            O => \N__45333\,
            I => \N__45294\
        );

    \I__10261\ : CascadeMux
    port map (
            O => \N__45332\,
            I => \N__45291\
        );

    \I__10260\ : InMux
    port map (
            O => \N__45329\,
            I => \N__45287\
        );

    \I__10259\ : InMux
    port map (
            O => \N__45326\,
            I => \N__45284\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__45323\,
            I => \N__45281\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__45320\,
            I => \N__45276\
        );

    \I__10256\ : Span4Mux_h
    port map (
            O => \N__45317\,
            I => \N__45276\
        );

    \I__10255\ : InMux
    port map (
            O => \N__45316\,
            I => \N__45271\
        );

    \I__10254\ : InMux
    port map (
            O => \N__45315\,
            I => \N__45271\
        );

    \I__10253\ : InMux
    port map (
            O => \N__45314\,
            I => \N__45268\
        );

    \I__10252\ : InMux
    port map (
            O => \N__45313\,
            I => \N__45265\
        );

    \I__10251\ : InMux
    port map (
            O => \N__45312\,
            I => \N__45260\
        );

    \I__10250\ : InMux
    port map (
            O => \N__45311\,
            I => \N__45260\
        );

    \I__10249\ : Span4Mux_v
    port map (
            O => \N__45306\,
            I => \N__45257\
        );

    \I__10248\ : InMux
    port map (
            O => \N__45303\,
            I => \N__45252\
        );

    \I__10247\ : InMux
    port map (
            O => \N__45300\,
            I => \N__45252\
        );

    \I__10246\ : InMux
    port map (
            O => \N__45297\,
            I => \N__45249\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__45294\,
            I => \N__45246\
        );

    \I__10244\ : InMux
    port map (
            O => \N__45291\,
            I => \N__45243\
        );

    \I__10243\ : InMux
    port map (
            O => \N__45290\,
            I => \N__45240\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__45287\,
            I => \N__45223\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__45284\,
            I => \N__45223\
        );

    \I__10240\ : Span12Mux_s11_v
    port map (
            O => \N__45281\,
            I => \N__45223\
        );

    \I__10239\ : Sp12to4
    port map (
            O => \N__45276\,
            I => \N__45223\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__45271\,
            I => \N__45223\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__45268\,
            I => \N__45223\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__45265\,
            I => \N__45223\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__45260\,
            I => \N__45223\
        );

    \I__10234\ : Odrv4
    port map (
            O => \N__45257\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__45252\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__45249\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10231\ : Odrv4
    port map (
            O => \N__45246\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__45243\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__45240\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10228\ : Odrv12
    port map (
            O => \N__45223\,
            I => \delay_measurement_inst.delay_tr9\
        );

    \I__10227\ : InMux
    port map (
            O => \N__45208\,
            I => \N__45205\
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__45205\,
            I => \N__45202\
        );

    \I__10225\ : Span12Mux_v
    port map (
            O => \N__45202\,
            I => \N__45199\
        );

    \I__10224\ : Odrv12
    port map (
            O => \N__45199\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\
        );

    \I__10223\ : InMux
    port map (
            O => \N__45196\,
            I => \N__45193\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__45193\,
            I => \N__45190\
        );

    \I__10221\ : Odrv4
    port map (
            O => \N__45190\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__10220\ : CascadeMux
    port map (
            O => \N__45187\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__10219\ : InMux
    port map (
            O => \N__45184\,
            I => \N__45181\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__45181\,
            I => \N__45177\
        );

    \I__10217\ : InMux
    port map (
            O => \N__45180\,
            I => \N__45174\
        );

    \I__10216\ : Odrv4
    port map (
            O => \N__45177\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__45174\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__10214\ : InMux
    port map (
            O => \N__45169\,
            I => \N__45165\
        );

    \I__10213\ : InMux
    port map (
            O => \N__45168\,
            I => \N__45162\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__45165\,
            I => \N__45159\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45156\
        );

    \I__10210\ : Span4Mux_h
    port map (
            O => \N__45159\,
            I => \N__45151\
        );

    \I__10209\ : Span4Mux_h
    port map (
            O => \N__45156\,
            I => \N__45151\
        );

    \I__10208\ : Odrv4
    port map (
            O => \N__45151\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10207\ : InMux
    port map (
            O => \N__45148\,
            I => \N__45144\
        );

    \I__10206\ : InMux
    port map (
            O => \N__45147\,
            I => \N__45141\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__45144\,
            I => \N__45138\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__45141\,
            I => \N__45135\
        );

    \I__10203\ : Span4Mux_v
    port map (
            O => \N__45138\,
            I => \N__45130\
        );

    \I__10202\ : Span4Mux_v
    port map (
            O => \N__45135\,
            I => \N__45130\
        );

    \I__10201\ : Odrv4
    port map (
            O => \N__45130\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__10200\ : CascadeMux
    port map (
            O => \N__45127\,
            I => \N__45124\
        );

    \I__10199\ : InMux
    port map (
            O => \N__45124\,
            I => \N__45120\
        );

    \I__10198\ : InMux
    port map (
            O => \N__45123\,
            I => \N__45117\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__45120\,
            I => \N__45114\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__45117\,
            I => \N__45111\
        );

    \I__10195\ : Span4Mux_v
    port map (
            O => \N__45114\,
            I => \N__45108\
        );

    \I__10194\ : Span4Mux_v
    port map (
            O => \N__45111\,
            I => \N__45105\
        );

    \I__10193\ : Sp12to4
    port map (
            O => \N__45108\,
            I => \N__45102\
        );

    \I__10192\ : Odrv4
    port map (
            O => \N__45105\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__10191\ : Odrv12
    port map (
            O => \N__45102\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__10190\ : InMux
    port map (
            O => \N__45097\,
            I => \N__45093\
        );

    \I__10189\ : InMux
    port map (
            O => \N__45096\,
            I => \N__45090\
        );

    \I__10188\ : LocalMux
    port map (
            O => \N__45093\,
            I => \N__45087\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__45090\,
            I => \N__45084\
        );

    \I__10186\ : Span4Mux_h
    port map (
            O => \N__45087\,
            I => \N__45081\
        );

    \I__10185\ : Odrv4
    port map (
            O => \N__45084\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__10184\ : Odrv4
    port map (
            O => \N__45081\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__10183\ : InMux
    port map (
            O => \N__45076\,
            I => \N__45073\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__45073\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19\
        );

    \I__10181\ : InMux
    port map (
            O => \N__45070\,
            I => \N__45067\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__45067\,
            I => \N__45064\
        );

    \I__10179\ : Span4Mux_h
    port map (
            O => \N__45064\,
            I => \N__45061\
        );

    \I__10178\ : Odrv4
    port map (
            O => \N__45061\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17\
        );

    \I__10177\ : CascadeMux
    port map (
            O => \N__45058\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18_cascade_\
        );

    \I__10176\ : InMux
    port map (
            O => \N__45055\,
            I => \N__45052\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__45052\,
            I => \N__45049\
        );

    \I__10174\ : Span4Mux_v
    port map (
            O => \N__45049\,
            I => \N__45046\
        );

    \I__10173\ : Odrv4
    port map (
            O => \N__45046\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16\
        );

    \I__10172\ : InMux
    port map (
            O => \N__45043\,
            I => \N__45040\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__45040\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25\
        );

    \I__10170\ : InMux
    port map (
            O => \N__45037\,
            I => \N__45034\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__45034\,
            I => \N__45031\
        );

    \I__10168\ : Span4Mux_h
    port map (
            O => \N__45031\,
            I => \N__45028\
        );

    \I__10167\ : Odrv4
    port map (
            O => \N__45028\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df28\
        );

    \I__10166\ : InMux
    port map (
            O => \N__45025\,
            I => \N__45022\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__45022\,
            I => \N__45019\
        );

    \I__10164\ : Span4Mux_h
    port map (
            O => \N__45019\,
            I => \N__45016\
        );

    \I__10163\ : Odrv4
    port map (
            O => \N__45016\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df26\
        );

    \I__10162\ : InMux
    port map (
            O => \N__45013\,
            I => \N__45010\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__45010\,
            I => \N__45007\
        );

    \I__10160\ : Span4Mux_v
    port map (
            O => \N__45007\,
            I => \N__45003\
        );

    \I__10159\ : InMux
    port map (
            O => \N__45006\,
            I => \N__45000\
        );

    \I__10158\ : Odrv4
    port map (
            O => \N__45003\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__45000\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__10156\ : CascadeMux
    port map (
            O => \N__44995\,
            I => \N__44991\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44994\,
            I => \N__44988\
        );

    \I__10154\ : InMux
    port map (
            O => \N__44991\,
            I => \N__44984\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__44988\,
            I => \N__44981\
        );

    \I__10152\ : CascadeMux
    port map (
            O => \N__44987\,
            I => \N__44978\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__44984\,
            I => \N__44975\
        );

    \I__10150\ : Span4Mux_v
    port map (
            O => \N__44981\,
            I => \N__44972\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44978\,
            I => \N__44968\
        );

    \I__10148\ : Span4Mux_v
    port map (
            O => \N__44975\,
            I => \N__44963\
        );

    \I__10147\ : Span4Mux_h
    port map (
            O => \N__44972\,
            I => \N__44963\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44971\,
            I => \N__44960\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__44968\,
            I => \elapsed_time_ns_1_RNI5GT8E1_0_13\
        );

    \I__10144\ : Odrv4
    port map (
            O => \N__44963\,
            I => \elapsed_time_ns_1_RNI5GT8E1_0_13\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__44960\,
            I => \elapsed_time_ns_1_RNI5GT8E1_0_13\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44950\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__44950\,
            I => \N__44947\
        );

    \I__10140\ : Span4Mux_h
    port map (
            O => \N__44947\,
            I => \N__44944\
        );

    \I__10139\ : Odrv4
    port map (
            O => \N__44944\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\
        );

    \I__10138\ : CascadeMux
    port map (
            O => \N__44941\,
            I => \N__44937\
        );

    \I__10137\ : CascadeMux
    port map (
            O => \N__44940\,
            I => \N__44934\
        );

    \I__10136\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44930\
        );

    \I__10135\ : InMux
    port map (
            O => \N__44934\,
            I => \N__44927\
        );

    \I__10134\ : InMux
    port map (
            O => \N__44933\,
            I => \N__44924\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__44930\,
            I => \N__44919\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__44927\,
            I => \N__44919\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__44924\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10130\ : Odrv12
    port map (
            O => \N__44919\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10129\ : InMux
    port map (
            O => \N__44914\,
            I => \N__44911\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__44911\,
            I => \N__44908\
        );

    \I__10127\ : Span4Mux_h
    port map (
            O => \N__44908\,
            I => \N__44904\
        );

    \I__10126\ : InMux
    port map (
            O => \N__44907\,
            I => \N__44901\
        );

    \I__10125\ : Span4Mux_v
    port map (
            O => \N__44904\,
            I => \N__44898\
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__44901\,
            I => \N__44895\
        );

    \I__10123\ : Odrv4
    port map (
            O => \N__44898\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__10122\ : Odrv4
    port map (
            O => \N__44895\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__10121\ : InMux
    port map (
            O => \N__44890\,
            I => \bfn_17_14_0_\
        );

    \I__10120\ : CascadeMux
    port map (
            O => \N__44887\,
            I => \N__44884\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44884\,
            I => \N__44880\
        );

    \I__10118\ : CascadeMux
    port map (
            O => \N__44883\,
            I => \N__44877\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__44880\,
            I => \N__44873\
        );

    \I__10116\ : InMux
    port map (
            O => \N__44877\,
            I => \N__44870\
        );

    \I__10115\ : InMux
    port map (
            O => \N__44876\,
            I => \N__44867\
        );

    \I__10114\ : Sp12to4
    port map (
            O => \N__44873\,
            I => \N__44862\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__44870\,
            I => \N__44862\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__44867\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10111\ : Odrv12
    port map (
            O => \N__44862\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10110\ : CascadeMux
    port map (
            O => \N__44857\,
            I => \N__44854\
        );

    \I__10109\ : InMux
    port map (
            O => \N__44854\,
            I => \N__44850\
        );

    \I__10108\ : CascadeMux
    port map (
            O => \N__44853\,
            I => \N__44847\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__44850\,
            I => \N__44844\
        );

    \I__10106\ : InMux
    port map (
            O => \N__44847\,
            I => \N__44841\
        );

    \I__10105\ : Span4Mux_h
    port map (
            O => \N__44844\,
            I => \N__44838\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__44841\,
            I => \N__44835\
        );

    \I__10103\ : Span4Mux_v
    port map (
            O => \N__44838\,
            I => \N__44830\
        );

    \I__10102\ : Span4Mux_h
    port map (
            O => \N__44835\,
            I => \N__44830\
        );

    \I__10101\ : Odrv4
    port map (
            O => \N__44830\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10100\ : InMux
    port map (
            O => \N__44827\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__10099\ : InMux
    port map (
            O => \N__44824\,
            I => \N__44820\
        );

    \I__10098\ : InMux
    port map (
            O => \N__44823\,
            I => \N__44817\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__44820\,
            I => \N__44814\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44817\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__10095\ : Odrv12
    port map (
            O => \N__44814\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__10094\ : CascadeMux
    port map (
            O => \N__44809\,
            I => \N__44806\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44806\,
            I => \N__44801\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44805\,
            I => \N__44798\
        );

    \I__10091\ : InMux
    port map (
            O => \N__44804\,
            I => \N__44795\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__44801\,
            I => \N__44790\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44798\,
            I => \N__44790\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__44795\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__10087\ : Odrv12
    port map (
            O => \N__44790\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__10086\ : InMux
    port map (
            O => \N__44785\,
            I => \N__44781\
        );

    \I__10085\ : InMux
    port map (
            O => \N__44784\,
            I => \N__44778\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__44781\,
            I => \N__44775\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__44778\,
            I => \N__44772\
        );

    \I__10082\ : Span4Mux_v
    port map (
            O => \N__44775\,
            I => \N__44769\
        );

    \I__10081\ : Span4Mux_h
    port map (
            O => \N__44772\,
            I => \N__44766\
        );

    \I__10080\ : Odrv4
    port map (
            O => \N__44769\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__10079\ : Odrv4
    port map (
            O => \N__44766\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44761\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__10077\ : InMux
    port map (
            O => \N__44758\,
            I => \N__44753\
        );

    \I__10076\ : InMux
    port map (
            O => \N__44757\,
            I => \N__44748\
        );

    \I__10075\ : InMux
    port map (
            O => \N__44756\,
            I => \N__44748\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__44753\,
            I => \N__44743\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__44748\,
            I => \N__44743\
        );

    \I__10072\ : Odrv12
    port map (
            O => \N__44743\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__10071\ : CascadeMux
    port map (
            O => \N__44740\,
            I => \N__44737\
        );

    \I__10070\ : InMux
    port map (
            O => \N__44737\,
            I => \N__44733\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44736\,
            I => \N__44730\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__44733\,
            I => \N__44727\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__44730\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__10066\ : Odrv12
    port map (
            O => \N__44727\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__10065\ : InMux
    port map (
            O => \N__44722\,
            I => \N__44718\
        );

    \I__10064\ : InMux
    port map (
            O => \N__44721\,
            I => \N__44715\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__44718\,
            I => \N__44712\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__44715\,
            I => \N__44709\
        );

    \I__10061\ : Span4Mux_v
    port map (
            O => \N__44712\,
            I => \N__44704\
        );

    \I__10060\ : Span4Mux_h
    port map (
            O => \N__44709\,
            I => \N__44704\
        );

    \I__10059\ : Odrv4
    port map (
            O => \N__44704\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__10058\ : InMux
    port map (
            O => \N__44701\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__10057\ : InMux
    port map (
            O => \N__44698\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__10056\ : InMux
    port map (
            O => \N__44695\,
            I => \N__44687\
        );

    \I__10055\ : InMux
    port map (
            O => \N__44694\,
            I => \N__44687\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44693\,
            I => \N__44684\
        );

    \I__10053\ : CascadeMux
    port map (
            O => \N__44692\,
            I => \N__44681\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__44687\,
            I => \N__44677\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__44684\,
            I => \N__44674\
        );

    \I__10050\ : InMux
    port map (
            O => \N__44681\,
            I => \N__44671\
        );

    \I__10049\ : InMux
    port map (
            O => \N__44680\,
            I => \N__44668\
        );

    \I__10048\ : Span4Mux_h
    port map (
            O => \N__44677\,
            I => \N__44665\
        );

    \I__10047\ : Span4Mux_h
    port map (
            O => \N__44674\,
            I => \N__44657\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__44671\,
            I => \N__44657\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__44668\,
            I => \N__44657\
        );

    \I__10044\ : Span4Mux_v
    port map (
            O => \N__44665\,
            I => \N__44654\
        );

    \I__10043\ : InMux
    port map (
            O => \N__44664\,
            I => \N__44651\
        );

    \I__10042\ : Span4Mux_v
    port map (
            O => \N__44657\,
            I => \N__44648\
        );

    \I__10041\ : Odrv4
    port map (
            O => \N__44654\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__10040\ : LocalMux
    port map (
            O => \N__44651\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__10039\ : Odrv4
    port map (
            O => \N__44648\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__10038\ : InMux
    port map (
            O => \N__44641\,
            I => \N__44637\
        );

    \I__10037\ : CascadeMux
    port map (
            O => \N__44640\,
            I => \N__44634\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__44637\,
            I => \N__44631\
        );

    \I__10035\ : InMux
    port map (
            O => \N__44634\,
            I => \N__44628\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__44631\,
            I => \N__44625\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__44628\,
            I => \N__44619\
        );

    \I__10032\ : Span4Mux_v
    port map (
            O => \N__44625\,
            I => \N__44619\
        );

    \I__10031\ : InMux
    port map (
            O => \N__44624\,
            I => \N__44615\
        );

    \I__10030\ : Span4Mux_v
    port map (
            O => \N__44619\,
            I => \N__44612\
        );

    \I__10029\ : InMux
    port map (
            O => \N__44618\,
            I => \N__44609\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__44615\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__10027\ : Odrv4
    port map (
            O => \N__44612\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__44609\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__10025\ : InMux
    port map (
            O => \N__44602\,
            I => \N__44598\
        );

    \I__10024\ : InMux
    port map (
            O => \N__44601\,
            I => \N__44594\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__44598\,
            I => \N__44591\
        );

    \I__10022\ : InMux
    port map (
            O => \N__44597\,
            I => \N__44588\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__44594\,
            I => \N__44585\
        );

    \I__10020\ : Span4Mux_v
    port map (
            O => \N__44591\,
            I => \N__44582\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__44588\,
            I => \N__44579\
        );

    \I__10018\ : Span4Mux_v
    port map (
            O => \N__44585\,
            I => \N__44576\
        );

    \I__10017\ : Span4Mux_v
    port map (
            O => \N__44582\,
            I => \N__44573\
        );

    \I__10016\ : Span4Mux_v
    port map (
            O => \N__44579\,
            I => \N__44570\
        );

    \I__10015\ : Span4Mux_v
    port map (
            O => \N__44576\,
            I => \N__44567\
        );

    \I__10014\ : Span4Mux_v
    port map (
            O => \N__44573\,
            I => \N__44562\
        );

    \I__10013\ : Span4Mux_h
    port map (
            O => \N__44570\,
            I => \N__44562\
        );

    \I__10012\ : Odrv4
    port map (
            O => \N__44567\,
            I => \il_min_comp1_D2\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__44562\,
            I => \il_min_comp1_D2\
        );

    \I__10010\ : InMux
    port map (
            O => \N__44557\,
            I => \N__44554\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__44554\,
            I => \N__44549\
        );

    \I__10008\ : InMux
    port map (
            O => \N__44553\,
            I => \N__44546\
        );

    \I__10007\ : InMux
    port map (
            O => \N__44552\,
            I => \N__44543\
        );

    \I__10006\ : Span4Mux_v
    port map (
            O => \N__44549\,
            I => \N__44536\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__44546\,
            I => \N__44536\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__44543\,
            I => \N__44533\
        );

    \I__10003\ : InMux
    port map (
            O => \N__44542\,
            I => \N__44529\
        );

    \I__10002\ : InMux
    port map (
            O => \N__44541\,
            I => \N__44526\
        );

    \I__10001\ : Span4Mux_h
    port map (
            O => \N__44536\,
            I => \N__44523\
        );

    \I__10000\ : Span4Mux_h
    port map (
            O => \N__44533\,
            I => \N__44520\
        );

    \I__9999\ : InMux
    port map (
            O => \N__44532\,
            I => \N__44517\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__44529\,
            I => \N__44512\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__44526\,
            I => \N__44512\
        );

    \I__9996\ : Odrv4
    port map (
            O => \N__44523\,
            I => phase_controller_inst1_state_4
        );

    \I__9995\ : Odrv4
    port map (
            O => \N__44520\,
            I => phase_controller_inst1_state_4
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__44517\,
            I => phase_controller_inst1_state_4
        );

    \I__9993\ : Odrv12
    port map (
            O => \N__44512\,
            I => phase_controller_inst1_state_4
        );

    \I__9992\ : InMux
    port map (
            O => \N__44503\,
            I => \N__44500\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__44500\,
            I => \N__44497\
        );

    \I__9990\ : Span4Mux_h
    port map (
            O => \N__44497\,
            I => \N__44494\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__44494\,
            I => \N__44491\
        );

    \I__9988\ : Span4Mux_h
    port map (
            O => \N__44491\,
            I => \N__44487\
        );

    \I__9987\ : InMux
    port map (
            O => \N__44490\,
            I => \N__44484\
        );

    \I__9986\ : Odrv4
    port map (
            O => \N__44487\,
            I => \phase_controller_inst1.N_55\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__44484\,
            I => \phase_controller_inst1.N_55\
        );

    \I__9984\ : CascadeMux
    port map (
            O => \N__44479\,
            I => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0_cascade_\
        );

    \I__9983\ : CascadeMux
    port map (
            O => \N__44476\,
            I => \N__44472\
        );

    \I__9982\ : CascadeMux
    port map (
            O => \N__44475\,
            I => \N__44469\
        );

    \I__9981\ : InMux
    port map (
            O => \N__44472\,
            I => \N__44466\
        );

    \I__9980\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44463\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__44466\,
            I => \N__44457\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__44463\,
            I => \N__44457\
        );

    \I__9977\ : InMux
    port map (
            O => \N__44462\,
            I => \N__44454\
        );

    \I__9976\ : Span4Mux_v
    port map (
            O => \N__44457\,
            I => \N__44451\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__44454\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__9974\ : Odrv4
    port map (
            O => \N__44451\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__9973\ : InMux
    port map (
            O => \N__44446\,
            I => \bfn_17_13_0_\
        );

    \I__9972\ : CascadeMux
    port map (
            O => \N__44443\,
            I => \N__44440\
        );

    \I__9971\ : InMux
    port map (
            O => \N__44440\,
            I => \N__44437\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__44437\,
            I => \N__44432\
        );

    \I__9969\ : InMux
    port map (
            O => \N__44436\,
            I => \N__44429\
        );

    \I__9968\ : InMux
    port map (
            O => \N__44435\,
            I => \N__44426\
        );

    \I__9967\ : Sp12to4
    port map (
            O => \N__44432\,
            I => \N__44421\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__44429\,
            I => \N__44421\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__44426\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9964\ : Odrv12
    port map (
            O => \N__44421\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__9963\ : InMux
    port map (
            O => \N__44416\,
            I => \N__44413\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__44413\,
            I => \N__44410\
        );

    \I__9961\ : Span4Mux_v
    port map (
            O => \N__44410\,
            I => \N__44406\
        );

    \I__9960\ : InMux
    port map (
            O => \N__44409\,
            I => \N__44403\
        );

    \I__9959\ : Odrv4
    port map (
            O => \N__44406\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__44403\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9957\ : InMux
    port map (
            O => \N__44398\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__9956\ : InMux
    port map (
            O => \N__44395\,
            I => \N__44388\
        );

    \I__9955\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44388\
        );

    \I__9954\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44385\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__44388\,
            I => \N__44382\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__44385\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__9951\ : Odrv12
    port map (
            O => \N__44382\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__9950\ : InMux
    port map (
            O => \N__44377\,
            I => \N__44374\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__44374\,
            I => \N__44371\
        );

    \I__9948\ : Span4Mux_h
    port map (
            O => \N__44371\,
            I => \N__44367\
        );

    \I__9947\ : InMux
    port map (
            O => \N__44370\,
            I => \N__44364\
        );

    \I__9946\ : Odrv4
    port map (
            O => \N__44367\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__44364\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9944\ : InMux
    port map (
            O => \N__44359\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__9943\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44349\
        );

    \I__9942\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44349\
        );

    \I__9941\ : InMux
    port map (
            O => \N__44354\,
            I => \N__44346\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__44349\,
            I => \N__44343\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__44346\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__9938\ : Odrv12
    port map (
            O => \N__44343\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__9937\ : InMux
    port map (
            O => \N__44338\,
            I => \N__44335\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__44335\,
            I => \N__44332\
        );

    \I__9935\ : Span4Mux_h
    port map (
            O => \N__44332\,
            I => \N__44328\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44331\,
            I => \N__44325\
        );

    \I__9933\ : Odrv4
    port map (
            O => \N__44328\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__44325\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__9931\ : InMux
    port map (
            O => \N__44320\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__9930\ : CascadeMux
    port map (
            O => \N__44317\,
            I => \N__44313\
        );

    \I__9929\ : CascadeMux
    port map (
            O => \N__44316\,
            I => \N__44310\
        );

    \I__9928\ : InMux
    port map (
            O => \N__44313\,
            I => \N__44304\
        );

    \I__9927\ : InMux
    port map (
            O => \N__44310\,
            I => \N__44304\
        );

    \I__9926\ : InMux
    port map (
            O => \N__44309\,
            I => \N__44301\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__44304\,
            I => \N__44298\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__44301\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__9923\ : Odrv12
    port map (
            O => \N__44298\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__9922\ : InMux
    port map (
            O => \N__44293\,
            I => \N__44290\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__44290\,
            I => \N__44286\
        );

    \I__9920\ : InMux
    port map (
            O => \N__44289\,
            I => \N__44283\
        );

    \I__9919\ : Span4Mux_v
    port map (
            O => \N__44286\,
            I => \N__44278\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__44283\,
            I => \N__44278\
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__44278\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__9916\ : InMux
    port map (
            O => \N__44275\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__9915\ : CascadeMux
    port map (
            O => \N__44272\,
            I => \N__44268\
        );

    \I__9914\ : CascadeMux
    port map (
            O => \N__44271\,
            I => \N__44265\
        );

    \I__9913\ : InMux
    port map (
            O => \N__44268\,
            I => \N__44259\
        );

    \I__9912\ : InMux
    port map (
            O => \N__44265\,
            I => \N__44259\
        );

    \I__9911\ : InMux
    port map (
            O => \N__44264\,
            I => \N__44256\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__44259\,
            I => \N__44253\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__44256\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__9908\ : Odrv12
    port map (
            O => \N__44253\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__9907\ : InMux
    port map (
            O => \N__44248\,
            I => \N__44245\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__44245\,
            I => \N__44241\
        );

    \I__9905\ : InMux
    port map (
            O => \N__44244\,
            I => \N__44238\
        );

    \I__9904\ : Span4Mux_h
    port map (
            O => \N__44241\,
            I => \N__44233\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__44238\,
            I => \N__44233\
        );

    \I__9902\ : Odrv4
    port map (
            O => \N__44233\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__9901\ : InMux
    port map (
            O => \N__44230\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__9900\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44221\
        );

    \I__9899\ : InMux
    port map (
            O => \N__44226\,
            I => \N__44221\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__44221\,
            I => \N__44217\
        );

    \I__9897\ : InMux
    port map (
            O => \N__44220\,
            I => \N__44214\
        );

    \I__9896\ : Span4Mux_v
    port map (
            O => \N__44217\,
            I => \N__44211\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__44214\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__9894\ : Odrv4
    port map (
            O => \N__44211\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__9893\ : CascadeMux
    port map (
            O => \N__44206\,
            I => \N__44203\
        );

    \I__9892\ : InMux
    port map (
            O => \N__44203\,
            I => \N__44200\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__44200\,
            I => \N__44197\
        );

    \I__9890\ : Span12Mux_v
    port map (
            O => \N__44197\,
            I => \N__44193\
        );

    \I__9889\ : InMux
    port map (
            O => \N__44196\,
            I => \N__44190\
        );

    \I__9888\ : Odrv12
    port map (
            O => \N__44193\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__44190\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__9886\ : InMux
    port map (
            O => \N__44185\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__9885\ : InMux
    port map (
            O => \N__44182\,
            I => \N__44176\
        );

    \I__9884\ : InMux
    port map (
            O => \N__44181\,
            I => \N__44176\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__44176\,
            I => \N__44172\
        );

    \I__9882\ : InMux
    port map (
            O => \N__44175\,
            I => \N__44169\
        );

    \I__9881\ : Span4Mux_v
    port map (
            O => \N__44172\,
            I => \N__44166\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__44169\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9879\ : Odrv4
    port map (
            O => \N__44166\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__9878\ : InMux
    port map (
            O => \N__44161\,
            I => \N__44158\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__44158\,
            I => \N__44154\
        );

    \I__9876\ : InMux
    port map (
            O => \N__44157\,
            I => \N__44151\
        );

    \I__9875\ : Span4Mux_h
    port map (
            O => \N__44154\,
            I => \N__44148\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__44151\,
            I => \N__44145\
        );

    \I__9873\ : Span4Mux_v
    port map (
            O => \N__44148\,
            I => \N__44142\
        );

    \I__9872\ : Span4Mux_h
    port map (
            O => \N__44145\,
            I => \N__44139\
        );

    \I__9871\ : Odrv4
    port map (
            O => \N__44142\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9870\ : Odrv4
    port map (
            O => \N__44139\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__9869\ : InMux
    port map (
            O => \N__44134\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__9868\ : CascadeMux
    port map (
            O => \N__44131\,
            I => \N__44128\
        );

    \I__9867\ : InMux
    port map (
            O => \N__44128\,
            I => \N__44124\
        );

    \I__9866\ : CascadeMux
    port map (
            O => \N__44127\,
            I => \N__44121\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__44124\,
            I => \N__44117\
        );

    \I__9864\ : InMux
    port map (
            O => \N__44121\,
            I => \N__44114\
        );

    \I__9863\ : InMux
    port map (
            O => \N__44120\,
            I => \N__44111\
        );

    \I__9862\ : Sp12to4
    port map (
            O => \N__44117\,
            I => \N__44106\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__44114\,
            I => \N__44106\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__44111\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__9859\ : Odrv12
    port map (
            O => \N__44106\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__9858\ : InMux
    port map (
            O => \N__44101\,
            I => \N__44098\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__44098\,
            I => \N__44095\
        );

    \I__9856\ : Span4Mux_v
    port map (
            O => \N__44095\,
            I => \N__44091\
        );

    \I__9855\ : InMux
    port map (
            O => \N__44094\,
            I => \N__44088\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__44091\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__44088\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__9852\ : InMux
    port map (
            O => \N__44083\,
            I => \bfn_17_12_0_\
        );

    \I__9851\ : CascadeMux
    port map (
            O => \N__44080\,
            I => \N__44076\
        );

    \I__9850\ : CascadeMux
    port map (
            O => \N__44079\,
            I => \N__44073\
        );

    \I__9849\ : InMux
    port map (
            O => \N__44076\,
            I => \N__44069\
        );

    \I__9848\ : InMux
    port map (
            O => \N__44073\,
            I => \N__44066\
        );

    \I__9847\ : InMux
    port map (
            O => \N__44072\,
            I => \N__44063\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__44069\,
            I => \N__44058\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__44066\,
            I => \N__44058\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__44063\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__9843\ : Odrv12
    port map (
            O => \N__44058\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__9842\ : InMux
    port map (
            O => \N__44053\,
            I => \N__44050\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__44050\,
            I => \N__44047\
        );

    \I__9840\ : Span4Mux_h
    port map (
            O => \N__44047\,
            I => \N__44043\
        );

    \I__9839\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44040\
        );

    \I__9838\ : Odrv4
    port map (
            O => \N__44043\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__44040\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__9836\ : InMux
    port map (
            O => \N__44035\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__9835\ : InMux
    port map (
            O => \N__44032\,
            I => \N__44026\
        );

    \I__9834\ : InMux
    port map (
            O => \N__44031\,
            I => \N__44026\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__44026\,
            I => \N__44022\
        );

    \I__9832\ : InMux
    port map (
            O => \N__44025\,
            I => \N__44019\
        );

    \I__9831\ : Span4Mux_v
    port map (
            O => \N__44022\,
            I => \N__44016\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__44019\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__9829\ : Odrv4
    port map (
            O => \N__44016\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__9828\ : InMux
    port map (
            O => \N__44011\,
            I => \N__44008\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__44008\,
            I => \N__44004\
        );

    \I__9826\ : CascadeMux
    port map (
            O => \N__44007\,
            I => \N__44001\
        );

    \I__9825\ : Span4Mux_v
    port map (
            O => \N__44004\,
            I => \N__43998\
        );

    \I__9824\ : InMux
    port map (
            O => \N__44001\,
            I => \N__43995\
        );

    \I__9823\ : Odrv4
    port map (
            O => \N__43998\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9822\ : LocalMux
    port map (
            O => \N__43995\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43990\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__9820\ : CascadeMux
    port map (
            O => \N__43987\,
            I => \N__43984\
        );

    \I__9819\ : InMux
    port map (
            O => \N__43984\,
            I => \N__43981\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__43981\,
            I => \N__43977\
        );

    \I__9817\ : InMux
    port map (
            O => \N__43980\,
            I => \N__43974\
        );

    \I__9816\ : Span4Mux_h
    port map (
            O => \N__43977\,
            I => \N__43968\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__43974\,
            I => \N__43968\
        );

    \I__9814\ : InMux
    port map (
            O => \N__43973\,
            I => \N__43965\
        );

    \I__9813\ : Span4Mux_v
    port map (
            O => \N__43968\,
            I => \N__43962\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__43965\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__9811\ : Odrv4
    port map (
            O => \N__43962\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__9810\ : InMux
    port map (
            O => \N__43957\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__9809\ : CascadeMux
    port map (
            O => \N__43954\,
            I => \N__43950\
        );

    \I__9808\ : CascadeMux
    port map (
            O => \N__43953\,
            I => \N__43947\
        );

    \I__9807\ : InMux
    port map (
            O => \N__43950\,
            I => \N__43941\
        );

    \I__9806\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43941\
        );

    \I__9805\ : InMux
    port map (
            O => \N__43946\,
            I => \N__43938\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__43941\,
            I => \N__43935\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__43938\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__9802\ : Odrv12
    port map (
            O => \N__43935\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43930\,
            I => \N__43926\
        );

    \I__9800\ : InMux
    port map (
            O => \N__43929\,
            I => \N__43923\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__43926\,
            I => \N__43920\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__43923\,
            I => \N__43917\
        );

    \I__9797\ : Span4Mux_h
    port map (
            O => \N__43920\,
            I => \N__43911\
        );

    \I__9796\ : Span4Mux_v
    port map (
            O => \N__43917\,
            I => \N__43911\
        );

    \I__9795\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43908\
        );

    \I__9794\ : Odrv4
    port map (
            O => \N__43911\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__43908\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\
        );

    \I__9792\ : InMux
    port map (
            O => \N__43903\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__9791\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43893\
        );

    \I__9790\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43893\
        );

    \I__9789\ : InMux
    port map (
            O => \N__43898\,
            I => \N__43890\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__43893\,
            I => \N__43887\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__43890\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__9786\ : Odrv12
    port map (
            O => \N__43887\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__9785\ : InMux
    port map (
            O => \N__43882\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__9784\ : InMux
    port map (
            O => \N__43879\,
            I => \N__43873\
        );

    \I__9783\ : InMux
    port map (
            O => \N__43878\,
            I => \N__43873\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__43873\,
            I => \N__43869\
        );

    \I__9781\ : InMux
    port map (
            O => \N__43872\,
            I => \N__43866\
        );

    \I__9780\ : Span4Mux_v
    port map (
            O => \N__43869\,
            I => \N__43863\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__43866\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__9778\ : Odrv4
    port map (
            O => \N__43863\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__9777\ : InMux
    port map (
            O => \N__43858\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__9776\ : CascadeMux
    port map (
            O => \N__43855\,
            I => \N__43851\
        );

    \I__9775\ : CascadeMux
    port map (
            O => \N__43854\,
            I => \N__43848\
        );

    \I__9774\ : InMux
    port map (
            O => \N__43851\,
            I => \N__43843\
        );

    \I__9773\ : InMux
    port map (
            O => \N__43848\,
            I => \N__43843\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__43843\,
            I => \N__43839\
        );

    \I__9771\ : InMux
    port map (
            O => \N__43842\,
            I => \N__43836\
        );

    \I__9770\ : Span4Mux_v
    port map (
            O => \N__43839\,
            I => \N__43833\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__43836\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__9768\ : Odrv4
    port map (
            O => \N__43833\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__9767\ : InMux
    port map (
            O => \N__43828\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43799\
        );

    \I__9765\ : InMux
    port map (
            O => \N__43824\,
            I => \N__43799\
        );

    \I__9764\ : InMux
    port map (
            O => \N__43823\,
            I => \N__43799\
        );

    \I__9763\ : InMux
    port map (
            O => \N__43822\,
            I => \N__43799\
        );

    \I__9762\ : InMux
    port map (
            O => \N__43821\,
            I => \N__43790\
        );

    \I__9761\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43790\
        );

    \I__9760\ : InMux
    port map (
            O => \N__43819\,
            I => \N__43790\
        );

    \I__9759\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43790\
        );

    \I__9758\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43781\
        );

    \I__9757\ : InMux
    port map (
            O => \N__43816\,
            I => \N__43781\
        );

    \I__9756\ : InMux
    port map (
            O => \N__43815\,
            I => \N__43781\
        );

    \I__9755\ : InMux
    port map (
            O => \N__43814\,
            I => \N__43781\
        );

    \I__9754\ : InMux
    port map (
            O => \N__43813\,
            I => \N__43764\
        );

    \I__9753\ : InMux
    port map (
            O => \N__43812\,
            I => \N__43764\
        );

    \I__9752\ : InMux
    port map (
            O => \N__43811\,
            I => \N__43755\
        );

    \I__9751\ : InMux
    port map (
            O => \N__43810\,
            I => \N__43755\
        );

    \I__9750\ : InMux
    port map (
            O => \N__43809\,
            I => \N__43755\
        );

    \I__9749\ : InMux
    port map (
            O => \N__43808\,
            I => \N__43755\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__43799\,
            I => \N__43748\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__43790\,
            I => \N__43748\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__43781\,
            I => \N__43748\
        );

    \I__9745\ : InMux
    port map (
            O => \N__43780\,
            I => \N__43739\
        );

    \I__9744\ : InMux
    port map (
            O => \N__43779\,
            I => \N__43739\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43778\,
            I => \N__43739\
        );

    \I__9742\ : InMux
    port map (
            O => \N__43777\,
            I => \N__43739\
        );

    \I__9741\ : InMux
    port map (
            O => \N__43776\,
            I => \N__43730\
        );

    \I__9740\ : InMux
    port map (
            O => \N__43775\,
            I => \N__43730\
        );

    \I__9739\ : InMux
    port map (
            O => \N__43774\,
            I => \N__43730\
        );

    \I__9738\ : InMux
    port map (
            O => \N__43773\,
            I => \N__43730\
        );

    \I__9737\ : InMux
    port map (
            O => \N__43772\,
            I => \N__43721\
        );

    \I__9736\ : InMux
    port map (
            O => \N__43771\,
            I => \N__43721\
        );

    \I__9735\ : InMux
    port map (
            O => \N__43770\,
            I => \N__43721\
        );

    \I__9734\ : InMux
    port map (
            O => \N__43769\,
            I => \N__43721\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__43764\,
            I => \N__43718\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__43755\,
            I => \N__43715\
        );

    \I__9731\ : Span4Mux_v
    port map (
            O => \N__43748\,
            I => \N__43710\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__43739\,
            I => \N__43710\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__43730\,
            I => \N__43705\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__43721\,
            I => \N__43705\
        );

    \I__9727\ : Span4Mux_h
    port map (
            O => \N__43718\,
            I => \N__43700\
        );

    \I__9726\ : Span4Mux_h
    port map (
            O => \N__43715\,
            I => \N__43700\
        );

    \I__9725\ : Span4Mux_h
    port map (
            O => \N__43710\,
            I => \N__43697\
        );

    \I__9724\ : Odrv4
    port map (
            O => \N__43705\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9723\ : Odrv4
    port map (
            O => \N__43700\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9722\ : Odrv4
    port map (
            O => \N__43697\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9721\ : InMux
    port map (
            O => \N__43690\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__9720\ : CEMux
    port map (
            O => \N__43687\,
            I => \N__43684\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__43684\,
            I => \N__43680\
        );

    \I__9718\ : CEMux
    port map (
            O => \N__43683\,
            I => \N__43677\
        );

    \I__9717\ : Span4Mux_h
    port map (
            O => \N__43680\,
            I => \N__43670\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__43677\,
            I => \N__43670\
        );

    \I__9715\ : CEMux
    port map (
            O => \N__43676\,
            I => \N__43667\
        );

    \I__9714\ : CEMux
    port map (
            O => \N__43675\,
            I => \N__43664\
        );

    \I__9713\ : Span4Mux_v
    port map (
            O => \N__43670\,
            I => \N__43661\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__43667\,
            I => \N__43658\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__43664\,
            I => \N__43655\
        );

    \I__9710\ : Span4Mux_h
    port map (
            O => \N__43661\,
            I => \N__43652\
        );

    \I__9709\ : Span4Mux_h
    port map (
            O => \N__43658\,
            I => \N__43649\
        );

    \I__9708\ : Span4Mux_h
    port map (
            O => \N__43655\,
            I => \N__43646\
        );

    \I__9707\ : Span4Mux_h
    port map (
            O => \N__43652\,
            I => \N__43643\
        );

    \I__9706\ : Span4Mux_h
    port map (
            O => \N__43649\,
            I => \N__43640\
        );

    \I__9705\ : Span4Mux_h
    port map (
            O => \N__43646\,
            I => \N__43637\
        );

    \I__9704\ : Odrv4
    port map (
            O => \N__43643\,
            I => \delay_measurement_inst.delay_tr_timer.N_400_i\
        );

    \I__9703\ : Odrv4
    port map (
            O => \N__43640\,
            I => \delay_measurement_inst.delay_tr_timer.N_400_i\
        );

    \I__9702\ : Odrv4
    port map (
            O => \N__43637\,
            I => \delay_measurement_inst.delay_tr_timer.N_400_i\
        );

    \I__9701\ : InMux
    port map (
            O => \N__43630\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__9700\ : InMux
    port map (
            O => \N__43627\,
            I => \N__43621\
        );

    \I__9699\ : InMux
    port map (
            O => \N__43626\,
            I => \N__43621\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__43621\,
            I => \N__43617\
        );

    \I__9697\ : InMux
    port map (
            O => \N__43620\,
            I => \N__43614\
        );

    \I__9696\ : Span4Mux_v
    port map (
            O => \N__43617\,
            I => \N__43611\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__43614\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__9694\ : Odrv4
    port map (
            O => \N__43611\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__9693\ : InMux
    port map (
            O => \N__43606\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__9692\ : InMux
    port map (
            O => \N__43603\,
            I => \N__43597\
        );

    \I__9691\ : InMux
    port map (
            O => \N__43602\,
            I => \N__43597\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__43597\,
            I => \N__43593\
        );

    \I__9689\ : InMux
    port map (
            O => \N__43596\,
            I => \N__43590\
        );

    \I__9688\ : Span4Mux_v
    port map (
            O => \N__43593\,
            I => \N__43587\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__43590\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__9686\ : Odrv4
    port map (
            O => \N__43587\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__9685\ : InMux
    port map (
            O => \N__43582\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__9684\ : CascadeMux
    port map (
            O => \N__43579\,
            I => \N__43575\
        );

    \I__9683\ : CascadeMux
    port map (
            O => \N__43578\,
            I => \N__43572\
        );

    \I__9682\ : InMux
    port map (
            O => \N__43575\,
            I => \N__43566\
        );

    \I__9681\ : InMux
    port map (
            O => \N__43572\,
            I => \N__43566\
        );

    \I__9680\ : InMux
    port map (
            O => \N__43571\,
            I => \N__43563\
        );

    \I__9679\ : LocalMux
    port map (
            O => \N__43566\,
            I => \N__43560\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__43563\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__9677\ : Odrv12
    port map (
            O => \N__43560\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__9676\ : InMux
    port map (
            O => \N__43555\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__9675\ : CascadeMux
    port map (
            O => \N__43552\,
            I => \N__43548\
        );

    \I__9674\ : CascadeMux
    port map (
            O => \N__43551\,
            I => \N__43545\
        );

    \I__9673\ : InMux
    port map (
            O => \N__43548\,
            I => \N__43539\
        );

    \I__9672\ : InMux
    port map (
            O => \N__43545\,
            I => \N__43539\
        );

    \I__9671\ : InMux
    port map (
            O => \N__43544\,
            I => \N__43536\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__43539\,
            I => \N__43533\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__43536\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__9668\ : Odrv12
    port map (
            O => \N__43533\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__9667\ : InMux
    port map (
            O => \N__43528\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__9666\ : InMux
    port map (
            O => \N__43525\,
            I => \N__43519\
        );

    \I__9665\ : InMux
    port map (
            O => \N__43524\,
            I => \N__43519\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__43519\,
            I => \N__43515\
        );

    \I__9663\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43512\
        );

    \I__9662\ : Span4Mux_v
    port map (
            O => \N__43515\,
            I => \N__43509\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__43512\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__9660\ : Odrv4
    port map (
            O => \N__43509\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__9659\ : InMux
    port map (
            O => \N__43504\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__9658\ : InMux
    port map (
            O => \N__43501\,
            I => \N__43495\
        );

    \I__9657\ : InMux
    port map (
            O => \N__43500\,
            I => \N__43495\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__43495\,
            I => \N__43491\
        );

    \I__9655\ : InMux
    port map (
            O => \N__43494\,
            I => \N__43488\
        );

    \I__9654\ : Span4Mux_v
    port map (
            O => \N__43491\,
            I => \N__43485\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__43488\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__9652\ : Odrv4
    port map (
            O => \N__43485\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__9651\ : InMux
    port map (
            O => \N__43480\,
            I => \N__43477\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__43477\,
            I => \N__43473\
        );

    \I__9649\ : InMux
    port map (
            O => \N__43476\,
            I => \N__43470\
        );

    \I__9648\ : Odrv12
    port map (
            O => \N__43473\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__43470\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9646\ : InMux
    port map (
            O => \N__43465\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__9645\ : InMux
    port map (
            O => \N__43462\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__9644\ : InMux
    port map (
            O => \N__43459\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__9643\ : InMux
    port map (
            O => \N__43456\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__9642\ : InMux
    port map (
            O => \N__43453\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__9641\ : InMux
    port map (
            O => \N__43450\,
            I => \bfn_17_10_0_\
        );

    \I__9640\ : InMux
    port map (
            O => \N__43447\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__9639\ : InMux
    port map (
            O => \N__43444\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__9638\ : InMux
    port map (
            O => \N__43441\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__9637\ : InMux
    port map (
            O => \N__43438\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__9636\ : InMux
    port map (
            O => \N__43435\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__9635\ : InMux
    port map (
            O => \N__43432\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__9634\ : InMux
    port map (
            O => \N__43429\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__9633\ : InMux
    port map (
            O => \N__43426\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__9632\ : InMux
    port map (
            O => \N__43423\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__9631\ : InMux
    port map (
            O => \N__43420\,
            I => \bfn_17_9_0_\
        );

    \I__9630\ : InMux
    port map (
            O => \N__43417\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__9629\ : InMux
    port map (
            O => \N__43414\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__9628\ : InMux
    port map (
            O => \N__43411\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__9627\ : InMux
    port map (
            O => \N__43408\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__9626\ : InMux
    port map (
            O => \N__43405\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__9625\ : InMux
    port map (
            O => \N__43402\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__9624\ : InMux
    port map (
            O => \N__43399\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__9623\ : InMux
    port map (
            O => \N__43396\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__9622\ : InMux
    port map (
            O => \N__43393\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__9621\ : InMux
    port map (
            O => \N__43390\,
            I => \bfn_17_8_0_\
        );

    \I__9620\ : InMux
    port map (
            O => \N__43387\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__9619\ : InMux
    port map (
            O => \N__43384\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__9618\ : CascadeMux
    port map (
            O => \N__43381\,
            I => \N__43378\
        );

    \I__9617\ : InMux
    port map (
            O => \N__43378\,
            I => \N__43372\
        );

    \I__9616\ : InMux
    port map (
            O => \N__43377\,
            I => \N__43369\
        );

    \I__9615\ : CascadeMux
    port map (
            O => \N__43376\,
            I => \N__43366\
        );

    \I__9614\ : InMux
    port map (
            O => \N__43375\,
            I => \N__43363\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__43372\,
            I => \N__43358\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__43369\,
            I => \N__43358\
        );

    \I__9611\ : InMux
    port map (
            O => \N__43366\,
            I => \N__43355\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__43363\,
            I => \N__43352\
        );

    \I__9609\ : Odrv12
    port map (
            O => \N__43358\,
            I => \elapsed_time_ns_1_RNIHHC6P1_0_18\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__43355\,
            I => \elapsed_time_ns_1_RNIHHC6P1_0_18\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__43352\,
            I => \elapsed_time_ns_1_RNIHHC6P1_0_18\
        );

    \I__9606\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43341\
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__43344\,
            I => \N__43338\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__43341\,
            I => \N__43335\
        );

    \I__9603\ : InMux
    port map (
            O => \N__43338\,
            I => \N__43332\
        );

    \I__9602\ : Span12Mux_s8_v
    port map (
            O => \N__43335\,
            I => \N__43329\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__43332\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__9600\ : Odrv12
    port map (
            O => \N__43329\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__9599\ : InMux
    port map (
            O => \N__43324\,
            I => \N__43321\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__43321\,
            I => \N__43318\
        );

    \I__9597\ : Span4Mux_h
    port map (
            O => \N__43318\,
            I => \N__43315\
        );

    \I__9596\ : Span4Mux_h
    port map (
            O => \N__43315\,
            I => \N__43312\
        );

    \I__9595\ : Odrv4
    port map (
            O => \N__43312\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__9594\ : CascadeMux
    port map (
            O => \N__43309\,
            I => \N__43305\
        );

    \I__9593\ : InMux
    port map (
            O => \N__43308\,
            I => \N__43302\
        );

    \I__9592\ : InMux
    port map (
            O => \N__43305\,
            I => \N__43299\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__43302\,
            I => \N__43292\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__43299\,
            I => \N__43292\
        );

    \I__9589\ : InMux
    port map (
            O => \N__43298\,
            I => \N__43289\
        );

    \I__9588\ : InMux
    port map (
            O => \N__43297\,
            I => \N__43286\
        );

    \I__9587\ : Span4Mux_v
    port map (
            O => \N__43292\,
            I => \N__43281\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__43289\,
            I => \N__43281\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__43286\,
            I => \elapsed_time_ns_1_RNI2DT8E1_0_10\
        );

    \I__9584\ : Odrv4
    port map (
            O => \N__43281\,
            I => \elapsed_time_ns_1_RNI2DT8E1_0_10\
        );

    \I__9583\ : InMux
    port map (
            O => \N__43276\,
            I => \N__43273\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__43273\,
            I => \N__43270\
        );

    \I__9581\ : Span12Mux_h
    port map (
            O => \N__43270\,
            I => \N__43267\
        );

    \I__9580\ : Odrv12
    port map (
            O => \N__43267\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__9579\ : CascadeMux
    port map (
            O => \N__43264\,
            I => \N__43260\
        );

    \I__9578\ : InMux
    port map (
            O => \N__43263\,
            I => \N__43256\
        );

    \I__9577\ : InMux
    port map (
            O => \N__43260\,
            I => \N__43253\
        );

    \I__9576\ : CascadeMux
    port map (
            O => \N__43259\,
            I => \N__43250\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__43256\,
            I => \N__43244\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__43253\,
            I => \N__43244\
        );

    \I__9573\ : InMux
    port map (
            O => \N__43250\,
            I => \N__43239\
        );

    \I__9572\ : InMux
    port map (
            O => \N__43249\,
            I => \N__43239\
        );

    \I__9571\ : Odrv12
    port map (
            O => \N__43244\,
            I => \elapsed_time_ns_1_RNI3ET8E1_0_11\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__43239\,
            I => \elapsed_time_ns_1_RNI3ET8E1_0_11\
        );

    \I__9569\ : InMux
    port map (
            O => \N__43234\,
            I => \N__43231\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__43231\,
            I => \N__43228\
        );

    \I__9567\ : Span4Mux_h
    port map (
            O => \N__43228\,
            I => \N__43225\
        );

    \I__9566\ : Span4Mux_h
    port map (
            O => \N__43225\,
            I => \N__43222\
        );

    \I__9565\ : Odrv4
    port map (
            O => \N__43222\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__9564\ : CascadeMux
    port map (
            O => \N__43219\,
            I => \N__43216\
        );

    \I__9563\ : InMux
    port map (
            O => \N__43216\,
            I => \N__43212\
        );

    \I__9562\ : InMux
    port map (
            O => \N__43215\,
            I => \N__43209\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__43212\,
            I => \N__43203\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__43209\,
            I => \N__43203\
        );

    \I__9559\ : InMux
    port map (
            O => \N__43208\,
            I => \N__43200\
        );

    \I__9558\ : Odrv12
    port map (
            O => \N__43203\,
            I => \elapsed_time_ns_1_RNI4FT8E1_0_12\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__43200\,
            I => \elapsed_time_ns_1_RNI4FT8E1_0_12\
        );

    \I__9556\ : InMux
    port map (
            O => \N__43195\,
            I => \N__43192\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__43192\,
            I => \N__43189\
        );

    \I__9554\ : Span4Mux_h
    port map (
            O => \N__43189\,
            I => \N__43186\
        );

    \I__9553\ : Span4Mux_h
    port map (
            O => \N__43186\,
            I => \N__43183\
        );

    \I__9552\ : Odrv4
    port map (
            O => \N__43183\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__9551\ : InMux
    port map (
            O => \N__43180\,
            I => \N__43177\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__43177\,
            I => \N__43174\
        );

    \I__9549\ : Span4Mux_h
    port map (
            O => \N__43174\,
            I => \N__43171\
        );

    \I__9548\ : Span4Mux_h
    port map (
            O => \N__43171\,
            I => \N__43168\
        );

    \I__9547\ : Odrv4
    port map (
            O => \N__43168\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__9546\ : InMux
    port map (
            O => \N__43165\,
            I => \N__43162\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__43162\,
            I => \N__43159\
        );

    \I__9544\ : Span4Mux_h
    port map (
            O => \N__43159\,
            I => \N__43156\
        );

    \I__9543\ : Span4Mux_h
    port map (
            O => \N__43156\,
            I => \N__43153\
        );

    \I__9542\ : Odrv4
    port map (
            O => \N__43153\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__9541\ : CEMux
    port map (
            O => \N__43150\,
            I => \N__43145\
        );

    \I__9540\ : CEMux
    port map (
            O => \N__43149\,
            I => \N__43118\
        );

    \I__9539\ : CEMux
    port map (
            O => \N__43148\,
            I => \N__43115\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__43145\,
            I => \N__43112\
        );

    \I__9537\ : CEMux
    port map (
            O => \N__43144\,
            I => \N__43109\
        );

    \I__9536\ : CEMux
    port map (
            O => \N__43143\,
            I => \N__43106\
        );

    \I__9535\ : InMux
    port map (
            O => \N__43142\,
            I => \N__43097\
        );

    \I__9534\ : InMux
    port map (
            O => \N__43141\,
            I => \N__43097\
        );

    \I__9533\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43097\
        );

    \I__9532\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43097\
        );

    \I__9531\ : InMux
    port map (
            O => \N__43138\,
            I => \N__43082\
        );

    \I__9530\ : InMux
    port map (
            O => \N__43137\,
            I => \N__43082\
        );

    \I__9529\ : InMux
    port map (
            O => \N__43136\,
            I => \N__43082\
        );

    \I__9528\ : InMux
    port map (
            O => \N__43135\,
            I => \N__43073\
        );

    \I__9527\ : InMux
    port map (
            O => \N__43134\,
            I => \N__43073\
        );

    \I__9526\ : InMux
    port map (
            O => \N__43133\,
            I => \N__43073\
        );

    \I__9525\ : InMux
    port map (
            O => \N__43132\,
            I => \N__43073\
        );

    \I__9524\ : InMux
    port map (
            O => \N__43131\,
            I => \N__43064\
        );

    \I__9523\ : InMux
    port map (
            O => \N__43130\,
            I => \N__43064\
        );

    \I__9522\ : InMux
    port map (
            O => \N__43129\,
            I => \N__43064\
        );

    \I__9521\ : InMux
    port map (
            O => \N__43128\,
            I => \N__43064\
        );

    \I__9520\ : InMux
    port map (
            O => \N__43127\,
            I => \N__43055\
        );

    \I__9519\ : InMux
    port map (
            O => \N__43126\,
            I => \N__43055\
        );

    \I__9518\ : InMux
    port map (
            O => \N__43125\,
            I => \N__43055\
        );

    \I__9517\ : InMux
    port map (
            O => \N__43124\,
            I => \N__43055\
        );

    \I__9516\ : InMux
    port map (
            O => \N__43123\,
            I => \N__43048\
        );

    \I__9515\ : InMux
    port map (
            O => \N__43122\,
            I => \N__43048\
        );

    \I__9514\ : InMux
    port map (
            O => \N__43121\,
            I => \N__43048\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__43118\,
            I => \N__43043\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__43115\,
            I => \N__43043\
        );

    \I__9511\ : Span4Mux_v
    port map (
            O => \N__43112\,
            I => \N__43037\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__43109\,
            I => \N__43037\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__43106\,
            I => \N__43034\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__43097\,
            I => \N__43031\
        );

    \I__9507\ : InMux
    port map (
            O => \N__43096\,
            I => \N__43022\
        );

    \I__9506\ : InMux
    port map (
            O => \N__43095\,
            I => \N__43022\
        );

    \I__9505\ : InMux
    port map (
            O => \N__43094\,
            I => \N__43022\
        );

    \I__9504\ : InMux
    port map (
            O => \N__43093\,
            I => \N__43022\
        );

    \I__9503\ : InMux
    port map (
            O => \N__43092\,
            I => \N__43013\
        );

    \I__9502\ : InMux
    port map (
            O => \N__43091\,
            I => \N__43013\
        );

    \I__9501\ : InMux
    port map (
            O => \N__43090\,
            I => \N__43013\
        );

    \I__9500\ : InMux
    port map (
            O => \N__43089\,
            I => \N__43013\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__43082\,
            I => \N__43006\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__43073\,
            I => \N__43006\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__43064\,
            I => \N__43006\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__43055\,
            I => \N__43001\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__43048\,
            I => \N__43001\
        );

    \I__9494\ : Span4Mux_v
    port map (
            O => \N__43043\,
            I => \N__42998\
        );

    \I__9493\ : InMux
    port map (
            O => \N__43042\,
            I => \N__42995\
        );

    \I__9492\ : Span4Mux_h
    port map (
            O => \N__43037\,
            I => \N__42992\
        );

    \I__9491\ : Span4Mux_v
    port map (
            O => \N__43034\,
            I => \N__42979\
        );

    \I__9490\ : Span4Mux_v
    port map (
            O => \N__43031\,
            I => \N__42979\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__43022\,
            I => \N__42979\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__43013\,
            I => \N__42979\
        );

    \I__9487\ : Span4Mux_v
    port map (
            O => \N__43006\,
            I => \N__42979\
        );

    \I__9486\ : Span4Mux_v
    port map (
            O => \N__43001\,
            I => \N__42979\
        );

    \I__9485\ : Odrv4
    port map (
            O => \N__42998\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__42995\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__9483\ : Odrv4
    port map (
            O => \N__42992\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__9482\ : Odrv4
    port map (
            O => \N__42979\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__9481\ : InMux
    port map (
            O => \N__42970\,
            I => \bfn_17_7_0_\
        );

    \I__9480\ : InMux
    port map (
            O => \N__42967\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42964\,
            I => \N__42959\
        );

    \I__9478\ : InMux
    port map (
            O => \N__42963\,
            I => \N__42956\
        );

    \I__9477\ : InMux
    port map (
            O => \N__42962\,
            I => \N__42951\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__42959\,
            I => \N__42946\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__42956\,
            I => \N__42946\
        );

    \I__9474\ : InMux
    port map (
            O => \N__42955\,
            I => \N__42943\
        );

    \I__9473\ : InMux
    port map (
            O => \N__42954\,
            I => \N__42940\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__42951\,
            I => \elapsed_time_ns_1_RNIIIC6P1_0_19\
        );

    \I__9471\ : Odrv12
    port map (
            O => \N__42946\,
            I => \elapsed_time_ns_1_RNIIIC6P1_0_19\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__42943\,
            I => \elapsed_time_ns_1_RNIIIC6P1_0_19\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__42940\,
            I => \elapsed_time_ns_1_RNIIIC6P1_0_19\
        );

    \I__9468\ : CascadeMux
    port map (
            O => \N__42931\,
            I => \phase_controller_inst1.stoper_hc.N_318_cascade_\
        );

    \I__9467\ : InMux
    port map (
            O => \N__42928\,
            I => \N__42924\
        );

    \I__9466\ : InMux
    port map (
            O => \N__42927\,
            I => \N__42921\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__42924\,
            I => \N__42918\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__42921\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__9463\ : Odrv4
    port map (
            O => \N__42918\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__9462\ : InMux
    port map (
            O => \N__42913\,
            I => \N__42910\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__42910\,
            I => \N__42906\
        );

    \I__9460\ : InMux
    port map (
            O => \N__42909\,
            I => \N__42903\
        );

    \I__9459\ : Odrv4
    port map (
            O => \N__42906\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__42903\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__9457\ : InMux
    port map (
            O => \N__42898\,
            I => \N__42895\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__42895\,
            I => \N__42891\
        );

    \I__9455\ : InMux
    port map (
            O => \N__42894\,
            I => \N__42888\
        );

    \I__9454\ : Span4Mux_h
    port map (
            O => \N__42891\,
            I => \N__42885\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__42888\,
            I => \N__42882\
        );

    \I__9452\ : Span4Mux_v
    port map (
            O => \N__42885\,
            I => \N__42879\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__42882\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__9450\ : Odrv4
    port map (
            O => \N__42879\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__9449\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42871\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__42871\,
            I => \N__42867\
        );

    \I__9447\ : InMux
    port map (
            O => \N__42870\,
            I => \N__42863\
        );

    \I__9446\ : Span12Mux_v
    port map (
            O => \N__42867\,
            I => \N__42860\
        );

    \I__9445\ : InMux
    port map (
            O => \N__42866\,
            I => \N__42857\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__42863\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__9443\ : Odrv12
    port map (
            O => \N__42860\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__42857\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__9441\ : InMux
    port map (
            O => \N__42850\,
            I => \N__42847\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__42847\,
            I => \N__42843\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__42846\,
            I => \N__42839\
        );

    \I__9438\ : Span4Mux_h
    port map (
            O => \N__42843\,
            I => \N__42836\
        );

    \I__9437\ : InMux
    port map (
            O => \N__42842\,
            I => \N__42833\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42830\
        );

    \I__9435\ : Span4Mux_h
    port map (
            O => \N__42836\,
            I => \N__42827\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__42833\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__42830\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__42827\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__9431\ : CascadeMux
    port map (
            O => \N__42820\,
            I => \N__42817\
        );

    \I__9430\ : InMux
    port map (
            O => \N__42817\,
            I => \N__42814\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__42814\,
            I => \N__42811\
        );

    \I__9428\ : Span4Mux_h
    port map (
            O => \N__42811\,
            I => \N__42808\
        );

    \I__9427\ : Odrv4
    port map (
            O => \N__42808\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__9426\ : CascadeMux
    port map (
            O => \N__42805\,
            I => \N__42802\
        );

    \I__9425\ : InMux
    port map (
            O => \N__42802\,
            I => \N__42796\
        );

    \I__9424\ : InMux
    port map (
            O => \N__42801\,
            I => \N__42796\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__42796\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42793\,
            I => \N__42790\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__42790\,
            I => \N__42786\
        );

    \I__9420\ : InMux
    port map (
            O => \N__42789\,
            I => \N__42783\
        );

    \I__9419\ : Odrv4
    port map (
            O => \N__42786\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__42783\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__9417\ : CascadeMux
    port map (
            O => \N__42778\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_\
        );

    \I__9416\ : InMux
    port map (
            O => \N__42775\,
            I => \N__42770\
        );

    \I__9415\ : InMux
    port map (
            O => \N__42774\,
            I => \N__42766\
        );

    \I__9414\ : InMux
    port map (
            O => \N__42773\,
            I => \N__42763\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__42770\,
            I => \N__42760\
        );

    \I__9412\ : InMux
    port map (
            O => \N__42769\,
            I => \N__42757\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__42766\,
            I => \N__42752\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__42763\,
            I => \N__42752\
        );

    \I__9409\ : Span4Mux_v
    port map (
            O => \N__42760\,
            I => \N__42749\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__42757\,
            I => \elapsed_time_ns_1_RNIGGC6P1_0_17\
        );

    \I__9407\ : Odrv4
    port map (
            O => \N__42752\,
            I => \elapsed_time_ns_1_RNIGGC6P1_0_17\
        );

    \I__9406\ : Odrv4
    port map (
            O => \N__42749\,
            I => \elapsed_time_ns_1_RNIGGC6P1_0_17\
        );

    \I__9405\ : CascadeMux
    port map (
            O => \N__42742\,
            I => \elapsed_time_ns_1_RNIGGC6P1_0_17_cascade_\
        );

    \I__9404\ : CascadeMux
    port map (
            O => \N__42739\,
            I => \N__42736\
        );

    \I__9403\ : InMux
    port map (
            O => \N__42736\,
            I => \N__42733\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__42733\,
            I => \N__42730\
        );

    \I__9401\ : Span4Mux_v
    port map (
            O => \N__42730\,
            I => \N__42727\
        );

    \I__9400\ : Span4Mux_h
    port map (
            O => \N__42727\,
            I => \N__42724\
        );

    \I__9399\ : Odrv4
    port map (
            O => \N__42724\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__9398\ : CascadeMux
    port map (
            O => \N__42721\,
            I => \N__42718\
        );

    \I__9397\ : InMux
    port map (
            O => \N__42718\,
            I => \N__42712\
        );

    \I__9396\ : InMux
    port map (
            O => \N__42717\,
            I => \N__42712\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__42712\,
            I => \N__42709\
        );

    \I__9394\ : Span4Mux_h
    port map (
            O => \N__42709\,
            I => \N__42705\
        );

    \I__9393\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42702\
        );

    \I__9392\ : Span4Mux_h
    port map (
            O => \N__42705\,
            I => \N__42699\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__42702\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__9390\ : Odrv4
    port map (
            O => \N__42699\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__9389\ : CascadeMux
    port map (
            O => \N__42694\,
            I => \N__42691\
        );

    \I__9388\ : InMux
    port map (
            O => \N__42691\,
            I => \N__42685\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42690\,
            I => \N__42685\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__42685\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__9385\ : InMux
    port map (
            O => \N__42682\,
            I => \N__42676\
        );

    \I__9384\ : InMux
    port map (
            O => \N__42681\,
            I => \N__42676\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__42676\,
            I => \N__42672\
        );

    \I__9382\ : InMux
    port map (
            O => \N__42675\,
            I => \N__42669\
        );

    \I__9381\ : Span12Mux_h
    port map (
            O => \N__42672\,
            I => \N__42666\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__42669\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__9379\ : Odrv12
    port map (
            O => \N__42666\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__9378\ : InMux
    port map (
            O => \N__42661\,
            I => \N__42658\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__42658\,
            I => \N__42655\
        );

    \I__9376\ : Span4Mux_v
    port map (
            O => \N__42655\,
            I => \N__42652\
        );

    \I__9375\ : Span4Mux_h
    port map (
            O => \N__42652\,
            I => \N__42649\
        );

    \I__9374\ : Odrv4
    port map (
            O => \N__42649\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__9373\ : InMux
    port map (
            O => \N__42646\,
            I => \N__42640\
        );

    \I__9372\ : InMux
    port map (
            O => \N__42645\,
            I => \N__42637\
        );

    \I__9371\ : InMux
    port map (
            O => \N__42644\,
            I => \N__42634\
        );

    \I__9370\ : InMux
    port map (
            O => \N__42643\,
            I => \N__42631\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__42640\,
            I => \N__42628\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__42637\,
            I => \elapsed_time_ns_1_RNIFFC6P1_0_16\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__42634\,
            I => \elapsed_time_ns_1_RNIFFC6P1_0_16\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__42631\,
            I => \elapsed_time_ns_1_RNIFFC6P1_0_16\
        );

    \I__9365\ : Odrv4
    port map (
            O => \N__42628\,
            I => \elapsed_time_ns_1_RNIFFC6P1_0_16\
        );

    \I__9364\ : InMux
    port map (
            O => \N__42619\,
            I => \N__42613\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42618\,
            I => \N__42613\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__42613\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__9361\ : CascadeMux
    port map (
            O => \N__42610\,
            I => \N__42606\
        );

    \I__9360\ : InMux
    port map (
            O => \N__42609\,
            I => \N__42601\
        );

    \I__9359\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42601\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__42601\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__9357\ : InMux
    port map (
            O => \N__42598\,
            I => \N__42595\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__42595\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18\
        );

    \I__9355\ : CascadeMux
    port map (
            O => \N__42592\,
            I => \N__42588\
        );

    \I__9354\ : InMux
    port map (
            O => \N__42591\,
            I => \N__42583\
        );

    \I__9353\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42583\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__42583\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__9351\ : CascadeMux
    port map (
            O => \N__42580\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_\
        );

    \I__9350\ : InMux
    port map (
            O => \N__42577\,
            I => \N__42574\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__42574\,
            I => \N__42570\
        );

    \I__9348\ : InMux
    port map (
            O => \N__42573\,
            I => \N__42567\
        );

    \I__9347\ : Odrv4
    port map (
            O => \N__42570\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__42567\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__9345\ : CascadeMux
    port map (
            O => \N__42562\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\
        );

    \I__9344\ : CascadeMux
    port map (
            O => \N__42559\,
            I => \elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_\
        );

    \I__9343\ : InMux
    port map (
            O => \N__42556\,
            I => \N__42550\
        );

    \I__9342\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42550\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__42550\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__9340\ : InMux
    port map (
            O => \N__42547\,
            I => \N__42543\
        );

    \I__9339\ : InMux
    port map (
            O => \N__42546\,
            I => \N__42540\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__42543\,
            I => \N__42537\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__42540\,
            I => \N__42534\
        );

    \I__9336\ : Span4Mux_h
    port map (
            O => \N__42537\,
            I => \N__42531\
        );

    \I__9335\ : Odrv4
    port map (
            O => \N__42534\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9334\ : Odrv4
    port map (
            O => \N__42531\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9333\ : InMux
    port map (
            O => \N__42526\,
            I => \N__42522\
        );

    \I__9332\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42519\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__42522\,
            I => \N__42516\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__42519\,
            I => \N__42513\
        );

    \I__9329\ : Span4Mux_v
    port map (
            O => \N__42516\,
            I => \N__42508\
        );

    \I__9328\ : Span4Mux_h
    port map (
            O => \N__42513\,
            I => \N__42508\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__42508\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__9326\ : CascadeMux
    port map (
            O => \N__42505\,
            I => \N__42502\
        );

    \I__9325\ : InMux
    port map (
            O => \N__42502\,
            I => \N__42499\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__42499\,
            I => \elapsed_time_ns_1_RNIAMU8E1_0_27\
        );

    \I__9323\ : InMux
    port map (
            O => \N__42496\,
            I => \N__42490\
        );

    \I__9322\ : InMux
    port map (
            O => \N__42495\,
            I => \N__42490\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__42490\,
            I => \elapsed_time_ns_1_RNI9LU8E1_0_26\
        );

    \I__9320\ : InMux
    port map (
            O => \N__42487\,
            I => \N__42481\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42486\,
            I => \N__42481\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__42481\,
            I => \elapsed_time_ns_1_RNIBNU8E1_0_28\
        );

    \I__9317\ : CascadeMux
    port map (
            O => \N__42478\,
            I => \elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_\
        );

    \I__9316\ : CascadeMux
    port map (
            O => \N__42475\,
            I => \N__42472\
        );

    \I__9315\ : InMux
    port map (
            O => \N__42472\,
            I => \N__42468\
        );

    \I__9314\ : InMux
    port map (
            O => \N__42471\,
            I => \N__42465\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__42468\,
            I => \elapsed_time_ns_1_RNI8KU8E1_0_25\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__42465\,
            I => \elapsed_time_ns_1_RNI8KU8E1_0_25\
        );

    \I__9311\ : InMux
    port map (
            O => \N__42460\,
            I => \N__42457\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__42457\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15\
        );

    \I__9309\ : CascadeMux
    port map (
            O => \N__42454\,
            I => \N__42451\
        );

    \I__9308\ : InMux
    port map (
            O => \N__42451\,
            I => \N__42447\
        );

    \I__9307\ : InMux
    port map (
            O => \N__42450\,
            I => \N__42444\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__42447\,
            I => \elapsed_time_ns_1_RNI5HU8E1_0_22\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__42444\,
            I => \elapsed_time_ns_1_RNI5HU8E1_0_22\
        );

    \I__9304\ : CascadeMux
    port map (
            O => \N__42439\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15_cascade_\
        );

    \I__9303\ : CascadeMux
    port map (
            O => \N__42436\,
            I => \N__42433\
        );

    \I__9302\ : InMux
    port map (
            O => \N__42433\,
            I => \N__42429\
        );

    \I__9301\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42426\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__42429\,
            I => \elapsed_time_ns_1_RNI7JU8E1_0_24\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__42426\,
            I => \elapsed_time_ns_1_RNI7JU8E1_0_24\
        );

    \I__9298\ : CascadeMux
    port map (
            O => \N__42421\,
            I => \N__42418\
        );

    \I__9297\ : InMux
    port map (
            O => \N__42418\,
            I => \N__42414\
        );

    \I__9296\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42411\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__42414\,
            I => \elapsed_time_ns_1_RNI6IU8E1_0_23\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__42411\,
            I => \elapsed_time_ns_1_RNI6IU8E1_0_23\
        );

    \I__9293\ : InMux
    port map (
            O => \N__42406\,
            I => \N__42403\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__42403\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15\
        );

    \I__9291\ : InMux
    port map (
            O => \N__42400\,
            I => \N__42396\
        );

    \I__9290\ : InMux
    port map (
            O => \N__42399\,
            I => \N__42393\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__42396\,
            I => \N__42390\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__42393\,
            I => \N__42387\
        );

    \I__9287\ : Odrv4
    port map (
            O => \N__42390\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9286\ : Odrv4
    port map (
            O => \N__42387\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9285\ : InMux
    port map (
            O => \N__42382\,
            I => \N__42379\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__42379\,
            I => \N__42375\
        );

    \I__9283\ : InMux
    port map (
            O => \N__42378\,
            I => \N__42372\
        );

    \I__9282\ : Odrv4
    port map (
            O => \N__42375\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__42372\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__9280\ : InMux
    port map (
            O => \N__42367\,
            I => \N__42364\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__42364\,
            I => \N__42360\
        );

    \I__9278\ : InMux
    port map (
            O => \N__42363\,
            I => \N__42357\
        );

    \I__9277\ : Odrv4
    port map (
            O => \N__42360\,
            I => \delay_measurement_inst.delay_hc_timer.N_369\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__42357\,
            I => \delay_measurement_inst.delay_hc_timer.N_369\
        );

    \I__9275\ : CascadeMux
    port map (
            O => \N__42352\,
            I => \delay_measurement_inst.delay_hc_timer.N_344_i_cascade_\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__42349\,
            I => \elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_\
        );

    \I__9273\ : InMux
    port map (
            O => \N__42346\,
            I => \N__42340\
        );

    \I__9272\ : InMux
    port map (
            O => \N__42345\,
            I => \N__42340\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__42340\,
            I => \N__42337\
        );

    \I__9270\ : Span4Mux_h
    port map (
            O => \N__42337\,
            I => \N__42334\
        );

    \I__9269\ : Odrv4
    port map (
            O => \N__42334\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9268\ : InMux
    port map (
            O => \N__42331\,
            I => \N__42328\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__42328\,
            I => \N__42324\
        );

    \I__9266\ : InMux
    port map (
            O => \N__42327\,
            I => \N__42321\
        );

    \I__9265\ : Span4Mux_h
    port map (
            O => \N__42324\,
            I => \N__42318\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__42321\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__9263\ : Odrv4
    port map (
            O => \N__42318\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__9262\ : CascadeMux
    port map (
            O => \N__42313\,
            I => \N__42310\
        );

    \I__9261\ : InMux
    port map (
            O => \N__42310\,
            I => \N__42307\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__42307\,
            I => \N__42303\
        );

    \I__9259\ : InMux
    port map (
            O => \N__42306\,
            I => \N__42299\
        );

    \I__9258\ : Span4Mux_h
    port map (
            O => \N__42303\,
            I => \N__42296\
        );

    \I__9257\ : InMux
    port map (
            O => \N__42302\,
            I => \N__42293\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__42299\,
            I => \elapsed_time_ns_1_RNIMHKEE1_0_5\
        );

    \I__9255\ : Odrv4
    port map (
            O => \N__42296\,
            I => \elapsed_time_ns_1_RNIMHKEE1_0_5\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__42293\,
            I => \elapsed_time_ns_1_RNIMHKEE1_0_5\
        );

    \I__9253\ : InMux
    port map (
            O => \N__42286\,
            I => \N__42276\
        );

    \I__9252\ : CascadeMux
    port map (
            O => \N__42285\,
            I => \N__42273\
        );

    \I__9251\ : InMux
    port map (
            O => \N__42284\,
            I => \N__42268\
        );

    \I__9250\ : InMux
    port map (
            O => \N__42283\,
            I => \N__42256\
        );

    \I__9249\ : InMux
    port map (
            O => \N__42282\,
            I => \N__42256\
        );

    \I__9248\ : InMux
    port map (
            O => \N__42281\,
            I => \N__42256\
        );

    \I__9247\ : InMux
    port map (
            O => \N__42280\,
            I => \N__42256\
        );

    \I__9246\ : InMux
    port map (
            O => \N__42279\,
            I => \N__42256\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__42276\,
            I => \N__42253\
        );

    \I__9244\ : InMux
    port map (
            O => \N__42273\,
            I => \N__42248\
        );

    \I__9243\ : InMux
    port map (
            O => \N__42272\,
            I => \N__42248\
        );

    \I__9242\ : InMux
    port map (
            O => \N__42271\,
            I => \N__42245\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__42268\,
            I => \N__42242\
        );

    \I__9240\ : InMux
    port map (
            O => \N__42267\,
            I => \N__42239\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__42256\,
            I => \N__42228\
        );

    \I__9238\ : Span4Mux_h
    port map (
            O => \N__42253\,
            I => \N__42228\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__42248\,
            I => \N__42228\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__42245\,
            I => \N__42228\
        );

    \I__9235\ : Span4Mux_h
    port map (
            O => \N__42242\,
            I => \N__42228\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__42239\,
            I => \phase_controller_inst1.stoper_hc.N_330\
        );

    \I__9233\ : Odrv4
    port map (
            O => \N__42228\,
            I => \phase_controller_inst1.stoper_hc.N_330\
        );

    \I__9232\ : CascadeMux
    port map (
            O => \N__42223\,
            I => \elapsed_time_ns_1_RNIMHKEE1_0_5_cascade_\
        );

    \I__9231\ : CascadeMux
    port map (
            O => \N__42220\,
            I => \N__42217\
        );

    \I__9230\ : InMux
    port map (
            O => \N__42217\,
            I => \N__42209\
        );

    \I__9229\ : InMux
    port map (
            O => \N__42216\,
            I => \N__42206\
        );

    \I__9228\ : CascadeMux
    port map (
            O => \N__42215\,
            I => \N__42197\
        );

    \I__9227\ : CascadeMux
    port map (
            O => \N__42214\,
            I => \N__42194\
        );

    \I__9226\ : InMux
    port map (
            O => \N__42213\,
            I => \N__42189\
        );

    \I__9225\ : InMux
    port map (
            O => \N__42212\,
            I => \N__42186\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__42209\,
            I => \N__42181\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__42206\,
            I => \N__42181\
        );

    \I__9222\ : InMux
    port map (
            O => \N__42205\,
            I => \N__42178\
        );

    \I__9221\ : InMux
    port map (
            O => \N__42204\,
            I => \N__42173\
        );

    \I__9220\ : InMux
    port map (
            O => \N__42203\,
            I => \N__42173\
        );

    \I__9219\ : InMux
    port map (
            O => \N__42202\,
            I => \N__42162\
        );

    \I__9218\ : InMux
    port map (
            O => \N__42201\,
            I => \N__42162\
        );

    \I__9217\ : InMux
    port map (
            O => \N__42200\,
            I => \N__42162\
        );

    \I__9216\ : InMux
    port map (
            O => \N__42197\,
            I => \N__42162\
        );

    \I__9215\ : InMux
    port map (
            O => \N__42194\,
            I => \N__42162\
        );

    \I__9214\ : InMux
    port map (
            O => \N__42193\,
            I => \N__42157\
        );

    \I__9213\ : InMux
    port map (
            O => \N__42192\,
            I => \N__42157\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__42189\,
            I => \N__42154\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__42186\,
            I => \N__42149\
        );

    \I__9210\ : Span4Mux_h
    port map (
            O => \N__42181\,
            I => \N__42149\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__42178\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__42173\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__42162\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__42157\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__9205\ : Odrv4
    port map (
            O => \N__42154\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__9204\ : Odrv4
    port map (
            O => \N__42149\,
            I => \phase_controller_inst1.stoper_hc.N_328\
        );

    \I__9203\ : InMux
    port map (
            O => \N__42136\,
            I => \N__42132\
        );

    \I__9202\ : InMux
    port map (
            O => \N__42135\,
            I => \N__42129\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__42132\,
            I => \N__42124\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__42129\,
            I => \N__42124\
        );

    \I__9199\ : Span4Mux_v
    port map (
            O => \N__42124\,
            I => \N__42121\
        );

    \I__9198\ : Odrv4
    port map (
            O => \N__42121\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__9197\ : InMux
    port map (
            O => \N__42118\,
            I => \N__42114\
        );

    \I__9196\ : InMux
    port map (
            O => \N__42117\,
            I => \N__42111\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__42114\,
            I => \N__42106\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__42111\,
            I => \N__42106\
        );

    \I__9193\ : Odrv4
    port map (
            O => \N__42106\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__9192\ : CascadeMux
    port map (
            O => \N__42103\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19_cascade_\
        );

    \I__9191\ : CascadeMux
    port map (
            O => \N__42100\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_\
        );

    \I__9190\ : CascadeMux
    port map (
            O => \N__42097\,
            I => \elapsed_time_ns_1_RNI4FT8E1_0_12_cascade_\
        );

    \I__9189\ : InMux
    port map (
            O => \N__42094\,
            I => \N__42091\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__42091\,
            I => \N__42088\
        );

    \I__9187\ : Span4Mux_h
    port map (
            O => \N__42088\,
            I => \N__42085\
        );

    \I__9186\ : Odrv4
    port map (
            O => \N__42085\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15\
        );

    \I__9185\ : InMux
    port map (
            O => \N__42082\,
            I => \N__42079\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__42079\,
            I => \N__42076\
        );

    \I__9183\ : Span4Mux_h
    port map (
            O => \N__42076\,
            I => \N__42073\
        );

    \I__9182\ : Odrv4
    port map (
            O => \N__42073\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14\
        );

    \I__9181\ : CascadeMux
    port map (
            O => \N__42070\,
            I => \N__42067\
        );

    \I__9180\ : InMux
    port map (
            O => \N__42067\,
            I => \N__42064\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__42064\,
            I => \N__42061\
        );

    \I__9178\ : Span4Mux_h
    port map (
            O => \N__42061\,
            I => \N__42058\
        );

    \I__9177\ : Odrv4
    port map (
            O => \N__42058\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20\
        );

    \I__9176\ : CascadeMux
    port map (
            O => \N__42055\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_\
        );

    \I__9175\ : CascadeMux
    port map (
            O => \N__42052\,
            I => \delay_measurement_inst.delay_hc_timer.N_369_cascade_\
        );

    \I__9174\ : CascadeMux
    port map (
            O => \N__42049\,
            I => \delay_measurement_inst.delay_hc_timer.N_367_clk_cascade_\
        );

    \I__9173\ : InMux
    port map (
            O => \N__42046\,
            I => \N__42042\
        );

    \I__9172\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42039\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__42042\,
            I => \elapsed_time_ns_1_RNI3FU8E1_0_20\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__42039\,
            I => \elapsed_time_ns_1_RNI3FU8E1_0_20\
        );

    \I__9169\ : InMux
    port map (
            O => \N__42034\,
            I => \N__42030\
        );

    \I__9168\ : InMux
    port map (
            O => \N__42033\,
            I => \N__42027\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__42030\,
            I => \N__42024\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__42027\,
            I => \N__42021\
        );

    \I__9165\ : Odrv12
    port map (
            O => \N__42024\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__42021\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9163\ : CascadeMux
    port map (
            O => \N__42016\,
            I => \N__42012\
        );

    \I__9162\ : InMux
    port map (
            O => \N__42015\,
            I => \N__42009\
        );

    \I__9161\ : InMux
    port map (
            O => \N__42012\,
            I => \N__42006\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__42009\,
            I => \N__42003\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__42006\,
            I => \N__42000\
        );

    \I__9158\ : Span4Mux_v
    port map (
            O => \N__42003\,
            I => \N__41997\
        );

    \I__9157\ : Span4Mux_h
    port map (
            O => \N__42000\,
            I => \N__41994\
        );

    \I__9156\ : Odrv4
    port map (
            O => \N__41997\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9155\ : Odrv4
    port map (
            O => \N__41994\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9154\ : CascadeMux
    port map (
            O => \N__41989\,
            I => \N__41986\
        );

    \I__9153\ : InMux
    port map (
            O => \N__41986\,
            I => \N__41983\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__41983\,
            I => \N__41980\
        );

    \I__9151\ : Span4Mux_h
    port map (
            O => \N__41980\,
            I => \N__41977\
        );

    \I__9150\ : Odrv4
    port map (
            O => \N__41977\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41974\,
            I => \N__41971\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__41971\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__9147\ : InMux
    port map (
            O => \N__41968\,
            I => \N__41964\
        );

    \I__9146\ : InMux
    port map (
            O => \N__41967\,
            I => \N__41960\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__41964\,
            I => \N__41957\
        );

    \I__9144\ : InMux
    port map (
            O => \N__41963\,
            I => \N__41952\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__41960\,
            I => \N__41949\
        );

    \I__9142\ : Span4Mux_h
    port map (
            O => \N__41957\,
            I => \N__41946\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41956\,
            I => \N__41941\
        );

    \I__9140\ : InMux
    port map (
            O => \N__41955\,
            I => \N__41941\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__41952\,
            I => \elapsed_time_ns_1_RNI8765M1_0_16\
        );

    \I__9138\ : Odrv12
    port map (
            O => \N__41949\,
            I => \elapsed_time_ns_1_RNI8765M1_0_16\
        );

    \I__9137\ : Odrv4
    port map (
            O => \N__41946\,
            I => \elapsed_time_ns_1_RNI8765M1_0_16\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41941\,
            I => \elapsed_time_ns_1_RNI8765M1_0_16\
        );

    \I__9135\ : InMux
    port map (
            O => \N__41932\,
            I => \N__41926\
        );

    \I__9134\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41926\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__41926\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41923\,
            I => \N__41919\
        );

    \I__9131\ : InMux
    port map (
            O => \N__41922\,
            I => \N__41915\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__41919\,
            I => \N__41912\
        );

    \I__9129\ : CascadeMux
    port map (
            O => \N__41918\,
            I => \N__41908\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41915\,
            I => \N__41905\
        );

    \I__9127\ : Span4Mux_h
    port map (
            O => \N__41912\,
            I => \N__41902\
        );

    \I__9126\ : InMux
    port map (
            O => \N__41911\,
            I => \N__41899\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41908\,
            I => \N__41896\
        );

    \I__9124\ : Odrv4
    port map (
            O => \N__41905\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17\
        );

    \I__9123\ : Odrv4
    port map (
            O => \N__41902\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__41899\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__41896\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17\
        );

    \I__9120\ : CascadeMux
    port map (
            O => \N__41887\,
            I => \N__41884\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41884\,
            I => \N__41878\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41883\,
            I => \N__41878\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41878\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__9116\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41869\
        );

    \I__9115\ : InMux
    port map (
            O => \N__41874\,
            I => \N__41869\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__41869\,
            I => \N__41865\
        );

    \I__9113\ : InMux
    port map (
            O => \N__41868\,
            I => \N__41862\
        );

    \I__9112\ : Span4Mux_h
    port map (
            O => \N__41865\,
            I => \N__41857\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__41862\,
            I => \N__41854\
        );

    \I__9110\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41851\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41860\,
            I => \N__41848\
        );

    \I__9108\ : Odrv4
    port map (
            O => \N__41857\,
            I => \elapsed_time_ns_1_RNIBA65M1_0_19\
        );

    \I__9107\ : Odrv4
    port map (
            O => \N__41854\,
            I => \elapsed_time_ns_1_RNIBA65M1_0_19\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__41851\,
            I => \elapsed_time_ns_1_RNIBA65M1_0_19\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__41848\,
            I => \elapsed_time_ns_1_RNIBA65M1_0_19\
        );

    \I__9104\ : CascadeMux
    port map (
            O => \N__41839\,
            I => \N__41836\
        );

    \I__9103\ : InMux
    port map (
            O => \N__41836\,
            I => \N__41833\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__41833\,
            I => \N__41830\
        );

    \I__9101\ : Odrv4
    port map (
            O => \N__41830\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__9100\ : CascadeMux
    port map (
            O => \N__41827\,
            I => \N__41824\
        );

    \I__9099\ : InMux
    port map (
            O => \N__41824\,
            I => \N__41818\
        );

    \I__9098\ : InMux
    port map (
            O => \N__41823\,
            I => \N__41818\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__41818\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41812\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__41812\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__9094\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41787\
        );

    \I__9093\ : InMux
    port map (
            O => \N__41808\,
            I => \N__41787\
        );

    \I__9092\ : InMux
    port map (
            O => \N__41807\,
            I => \N__41787\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41787\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41787\
        );

    \I__9089\ : InMux
    port map (
            O => \N__41804\,
            I => \N__41782\
        );

    \I__9088\ : InMux
    port map (
            O => \N__41803\,
            I => \N__41782\
        );

    \I__9087\ : CascadeMux
    port map (
            O => \N__41802\,
            I => \N__41765\
        );

    \I__9086\ : InMux
    port map (
            O => \N__41801\,
            I => \N__41752\
        );

    \I__9085\ : InMux
    port map (
            O => \N__41800\,
            I => \N__41752\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41799\,
            I => \N__41752\
        );

    \I__9083\ : InMux
    port map (
            O => \N__41798\,
            I => \N__41752\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__41787\,
            I => \N__41746\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__41782\,
            I => \N__41743\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41781\,
            I => \N__41732\
        );

    \I__9079\ : InMux
    port map (
            O => \N__41780\,
            I => \N__41732\
        );

    \I__9078\ : InMux
    port map (
            O => \N__41779\,
            I => \N__41732\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41778\,
            I => \N__41732\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41777\,
            I => \N__41732\
        );

    \I__9075\ : InMux
    port map (
            O => \N__41776\,
            I => \N__41719\
        );

    \I__9074\ : InMux
    port map (
            O => \N__41775\,
            I => \N__41719\
        );

    \I__9073\ : InMux
    port map (
            O => \N__41774\,
            I => \N__41719\
        );

    \I__9072\ : InMux
    port map (
            O => \N__41773\,
            I => \N__41719\
        );

    \I__9071\ : InMux
    port map (
            O => \N__41772\,
            I => \N__41719\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41771\,
            I => \N__41719\
        );

    \I__9069\ : InMux
    port map (
            O => \N__41770\,
            I => \N__41716\
        );

    \I__9068\ : InMux
    port map (
            O => \N__41769\,
            I => \N__41707\
        );

    \I__9067\ : InMux
    port map (
            O => \N__41768\,
            I => \N__41707\
        );

    \I__9066\ : InMux
    port map (
            O => \N__41765\,
            I => \N__41707\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41707\
        );

    \I__9064\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41700\
        );

    \I__9063\ : InMux
    port map (
            O => \N__41762\,
            I => \N__41700\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41761\,
            I => \N__41700\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__41752\,
            I => \N__41695\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41751\,
            I => \N__41688\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41750\,
            I => \N__41688\
        );

    \I__9058\ : InMux
    port map (
            O => \N__41749\,
            I => \N__41688\
        );

    \I__9057\ : Span4Mux_v
    port map (
            O => \N__41746\,
            I => \N__41681\
        );

    \I__9056\ : Span4Mux_v
    port map (
            O => \N__41743\,
            I => \N__41681\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__41732\,
            I => \N__41681\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__41719\,
            I => \N__41672\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__41716\,
            I => \N__41672\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__41707\,
            I => \N__41672\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__41700\,
            I => \N__41672\
        );

    \I__9050\ : InMux
    port map (
            O => \N__41699\,
            I => \N__41667\
        );

    \I__9049\ : InMux
    port map (
            O => \N__41698\,
            I => \N__41667\
        );

    \I__9048\ : Odrv4
    port map (
            O => \N__41695\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__41688\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9046\ : Odrv4
    port map (
            O => \N__41681\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9045\ : Odrv4
    port map (
            O => \N__41672\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__41667\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31\
        );

    \I__9043\ : CascadeMux
    port map (
            O => \N__41656\,
            I => \N__41652\
        );

    \I__9042\ : CascadeMux
    port map (
            O => \N__41655\,
            I => \N__41649\
        );

    \I__9041\ : InMux
    port map (
            O => \N__41652\,
            I => \N__41638\
        );

    \I__9040\ : InMux
    port map (
            O => \N__41649\,
            I => \N__41638\
        );

    \I__9039\ : InMux
    port map (
            O => \N__41648\,
            I => \N__41638\
        );

    \I__9038\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41638\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__41638\,
            I => \N__41618\
        );

    \I__9036\ : InMux
    port map (
            O => \N__41637\,
            I => \N__41607\
        );

    \I__9035\ : InMux
    port map (
            O => \N__41636\,
            I => \N__41607\
        );

    \I__9034\ : InMux
    port map (
            O => \N__41635\,
            I => \N__41607\
        );

    \I__9033\ : InMux
    port map (
            O => \N__41634\,
            I => \N__41607\
        );

    \I__9032\ : InMux
    port map (
            O => \N__41633\,
            I => \N__41607\
        );

    \I__9031\ : CascadeMux
    port map (
            O => \N__41632\,
            I => \N__41604\
        );

    \I__9030\ : CascadeMux
    port map (
            O => \N__41631\,
            I => \N__41601\
        );

    \I__9029\ : CascadeMux
    port map (
            O => \N__41630\,
            I => \N__41597\
        );

    \I__9028\ : InMux
    port map (
            O => \N__41629\,
            I => \N__41586\
        );

    \I__9027\ : InMux
    port map (
            O => \N__41628\,
            I => \N__41586\
        );

    \I__9026\ : InMux
    port map (
            O => \N__41627\,
            I => \N__41586\
        );

    \I__9025\ : InMux
    port map (
            O => \N__41626\,
            I => \N__41583\
        );

    \I__9024\ : InMux
    port map (
            O => \N__41625\,
            I => \N__41578\
        );

    \I__9023\ : InMux
    port map (
            O => \N__41624\,
            I => \N__41578\
        );

    \I__9022\ : CascadeMux
    port map (
            O => \N__41623\,
            I => \N__41575\
        );

    \I__9021\ : CascadeMux
    port map (
            O => \N__41622\,
            I => \N__41572\
        );

    \I__9020\ : CascadeMux
    port map (
            O => \N__41621\,
            I => \N__41569\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__41618\,
            I => \N__41565\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__41607\,
            I => \N__41562\
        );

    \I__9017\ : InMux
    port map (
            O => \N__41604\,
            I => \N__41555\
        );

    \I__9016\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41555\
        );

    \I__9015\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41555\
        );

    \I__9014\ : InMux
    port map (
            O => \N__41597\,
            I => \N__41546\
        );

    \I__9013\ : InMux
    port map (
            O => \N__41596\,
            I => \N__41546\
        );

    \I__9012\ : InMux
    port map (
            O => \N__41595\,
            I => \N__41546\
        );

    \I__9011\ : InMux
    port map (
            O => \N__41594\,
            I => \N__41546\
        );

    \I__9010\ : InMux
    port map (
            O => \N__41593\,
            I => \N__41543\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__41586\,
            I => \N__41538\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__41583\,
            I => \N__41538\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__41578\,
            I => \N__41535\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41575\,
            I => \N__41526\
        );

    \I__9005\ : InMux
    port map (
            O => \N__41572\,
            I => \N__41526\
        );

    \I__9004\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41526\
        );

    \I__9003\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41526\
        );

    \I__9002\ : Span4Mux_v
    port map (
            O => \N__41565\,
            I => \N__41521\
        );

    \I__9001\ : Span4Mux_h
    port map (
            O => \N__41562\,
            I => \N__41521\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41555\,
            I => \N__41510\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__41546\,
            I => \N__41510\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__41543\,
            I => \N__41510\
        );

    \I__8997\ : Span4Mux_v
    port map (
            O => \N__41538\,
            I => \N__41510\
        );

    \I__8996\ : Span4Mux_h
    port map (
            O => \N__41535\,
            I => \N__41510\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__41526\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8994\ : Odrv4
    port map (
            O => \N__41521\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8993\ : Odrv4
    port map (
            O => \N__41510\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\
        );

    \I__8992\ : InMux
    port map (
            O => \N__41503\,
            I => \N__41499\
        );

    \I__8991\ : InMux
    port map (
            O => \N__41502\,
            I => \N__41495\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__41499\,
            I => \N__41492\
        );

    \I__8989\ : CascadeMux
    port map (
            O => \N__41498\,
            I => \N__41489\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__41495\,
            I => \N__41485\
        );

    \I__8987\ : Span4Mux_h
    port map (
            O => \N__41492\,
            I => \N__41482\
        );

    \I__8986\ : InMux
    port map (
            O => \N__41489\,
            I => \N__41479\
        );

    \I__8985\ : InMux
    port map (
            O => \N__41488\,
            I => \N__41476\
        );

    \I__8984\ : Odrv4
    port map (
            O => \N__41485\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18\
        );

    \I__8983\ : Odrv4
    port map (
            O => \N__41482\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__41479\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__41476\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18\
        );

    \I__8980\ : InMux
    port map (
            O => \N__41467\,
            I => \N__41461\
        );

    \I__8979\ : InMux
    port map (
            O => \N__41466\,
            I => \N__41461\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__41461\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__8977\ : InMux
    port map (
            O => \N__41458\,
            I => \N__41455\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__41455\,
            I => \N__41452\
        );

    \I__8975\ : Odrv4
    port map (
            O => \N__41452\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14\
        );

    \I__8974\ : CascadeMux
    port map (
            O => \N__41449\,
            I => \N__41445\
        );

    \I__8973\ : InMux
    port map (
            O => \N__41448\,
            I => \N__41440\
        );

    \I__8972\ : InMux
    port map (
            O => \N__41445\,
            I => \N__41437\
        );

    \I__8971\ : InMux
    port map (
            O => \N__41444\,
            I => \N__41434\
        );

    \I__8970\ : InMux
    port map (
            O => \N__41443\,
            I => \N__41429\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__41440\,
            I => \N__41426\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__41437\,
            I => \N__41421\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__41434\,
            I => \N__41421\
        );

    \I__8966\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41418\
        );

    \I__8965\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41415\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__41429\,
            I => \N__41412\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__41426\,
            I => \N__41409\
        );

    \I__8962\ : Span4Mux_v
    port map (
            O => \N__41421\,
            I => \N__41402\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__41418\,
            I => \N__41402\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__41415\,
            I => \N__41402\
        );

    \I__8959\ : Odrv12
    port map (
            O => \N__41412\,
            I => \elapsed_time_ns_1_RNI6565M1_0_14\
        );

    \I__8958\ : Odrv4
    port map (
            O => \N__41409\,
            I => \elapsed_time_ns_1_RNI6565M1_0_14\
        );

    \I__8957\ : Odrv4
    port map (
            O => \N__41402\,
            I => \elapsed_time_ns_1_RNI6565M1_0_14\
        );

    \I__8956\ : InMux
    port map (
            O => \N__41395\,
            I => \N__41392\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__41392\,
            I => \N__41388\
        );

    \I__8954\ : InMux
    port map (
            O => \N__41391\,
            I => \N__41385\
        );

    \I__8953\ : Odrv12
    port map (
            O => \N__41388\,
            I => \delay_measurement_inst.delay_tr_timer.N_395\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__41385\,
            I => \delay_measurement_inst.delay_tr_timer.N_395\
        );

    \I__8951\ : InMux
    port map (
            O => \N__41380\,
            I => \N__41377\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__41377\,
            I => \N__41373\
        );

    \I__8949\ : InMux
    port map (
            O => \N__41376\,
            I => \N__41370\
        );

    \I__8948\ : Odrv4
    port map (
            O => \N__41373\,
            I => \delay_measurement_inst.delay_tr_timer.N_375\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__41370\,
            I => \delay_measurement_inst.delay_tr_timer.N_375\
        );

    \I__8946\ : InMux
    port map (
            O => \N__41365\,
            I => \N__41355\
        );

    \I__8945\ : InMux
    port map (
            O => \N__41364\,
            I => \N__41348\
        );

    \I__8944\ : InMux
    port map (
            O => \N__41363\,
            I => \N__41348\
        );

    \I__8943\ : InMux
    port map (
            O => \N__41362\,
            I => \N__41348\
        );

    \I__8942\ : InMux
    port map (
            O => \N__41361\,
            I => \N__41339\
        );

    \I__8941\ : InMux
    port map (
            O => \N__41360\,
            I => \N__41339\
        );

    \I__8940\ : InMux
    port map (
            O => \N__41359\,
            I => \N__41339\
        );

    \I__8939\ : InMux
    port map (
            O => \N__41358\,
            I => \N__41339\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__41355\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__41348\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__41339\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\
        );

    \I__8935\ : InMux
    port map (
            O => \N__41332\,
            I => \N__41329\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__41329\,
            I => \N__41326\
        );

    \I__8933\ : Odrv4
    port map (
            O => \N__41326\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\
        );

    \I__8932\ : CascadeMux
    port map (
            O => \N__41323\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\
        );

    \I__8931\ : InMux
    port map (
            O => \N__41320\,
            I => \N__41312\
        );

    \I__8930\ : InMux
    port map (
            O => \N__41319\,
            I => \N__41312\
        );

    \I__8929\ : InMux
    port map (
            O => \N__41318\,
            I => \N__41307\
        );

    \I__8928\ : InMux
    port map (
            O => \N__41317\,
            I => \N__41304\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__41312\,
            I => \N__41301\
        );

    \I__8926\ : InMux
    port map (
            O => \N__41311\,
            I => \N__41296\
        );

    \I__8925\ : InMux
    port map (
            O => \N__41310\,
            I => \N__41296\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__41307\,
            I => \N__41291\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__41304\,
            I => \N__41291\
        );

    \I__8922\ : Span4Mux_v
    port map (
            O => \N__41301\,
            I => \N__41286\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__41296\,
            I => \N__41286\
        );

    \I__8920\ : Odrv4
    port map (
            O => \N__41291\,
            I => \elapsed_time_ns_1_RNIQENQL1_0_9\
        );

    \I__8919\ : Odrv4
    port map (
            O => \N__41286\,
            I => \elapsed_time_ns_1_RNIQENQL1_0_9\
        );

    \I__8918\ : CascadeMux
    port map (
            O => \N__41281\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_\
        );

    \I__8917\ : InMux
    port map (
            O => \N__41278\,
            I => \N__41275\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__41275\,
            I => \N__41271\
        );

    \I__8915\ : InMux
    port map (
            O => \N__41274\,
            I => \N__41268\
        );

    \I__8914\ : Odrv12
    port map (
            O => \N__41271\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__41268\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__8912\ : InMux
    port map (
            O => \N__41263\,
            I => \N__41256\
        );

    \I__8911\ : InMux
    port map (
            O => \N__41262\,
            I => \N__41256\
        );

    \I__8910\ : InMux
    port map (
            O => \N__41261\,
            I => \N__41253\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__41256\,
            I => \N__41250\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__41253\,
            I => \N__41247\
        );

    \I__8907\ : Span4Mux_h
    port map (
            O => \N__41250\,
            I => \N__41243\
        );

    \I__8906\ : Span4Mux_v
    port map (
            O => \N__41247\,
            I => \N__41240\
        );

    \I__8905\ : InMux
    port map (
            O => \N__41246\,
            I => \N__41237\
        );

    \I__8904\ : Span4Mux_v
    port map (
            O => \N__41243\,
            I => \N__41234\
        );

    \I__8903\ : Odrv4
    port map (
            O => \N__41240\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__41237\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__8901\ : Odrv4
    port map (
            O => \N__41234\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__8900\ : CascadeMux
    port map (
            O => \N__41227\,
            I => \N__41224\
        );

    \I__8899\ : InMux
    port map (
            O => \N__41224\,
            I => \N__41219\
        );

    \I__8898\ : InMux
    port map (
            O => \N__41223\,
            I => \N__41214\
        );

    \I__8897\ : InMux
    port map (
            O => \N__41222\,
            I => \N__41214\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__41219\,
            I => \N__41211\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__41214\,
            I => \N__41208\
        );

    \I__8894\ : Span12Mux_h
    port map (
            O => \N__41211\,
            I => \N__41205\
        );

    \I__8893\ : Span12Mux_v
    port map (
            O => \N__41208\,
            I => \N__41200\
        );

    \I__8892\ : Span12Mux_v
    port map (
            O => \N__41205\,
            I => \N__41200\
        );

    \I__8891\ : Odrv12
    port map (
            O => \N__41200\,
            I => \il_max_comp2_D2\
        );

    \I__8890\ : InMux
    port map (
            O => \N__41197\,
            I => \N__41194\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__41194\,
            I => \N__41191\
        );

    \I__8888\ : Span4Mux_h
    port map (
            O => \N__41191\,
            I => \N__41186\
        );

    \I__8887\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41181\
        );

    \I__8886\ : InMux
    port map (
            O => \N__41189\,
            I => \N__41181\
        );

    \I__8885\ : Odrv4
    port map (
            O => \N__41186\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__41181\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__8883\ : CascadeMux
    port map (
            O => \N__41176\,
            I => \delay_measurement_inst.delay_tr_timer.N_353_cascade_\
        );

    \I__8882\ : InMux
    port map (
            O => \N__41173\,
            I => \N__41170\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__41170\,
            I => \N__41165\
        );

    \I__8880\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41160\
        );

    \I__8879\ : InMux
    port map (
            O => \N__41168\,
            I => \N__41160\
        );

    \I__8878\ : Odrv4
    port map (
            O => \N__41165\,
            I => \delay_measurement_inst.delay_tr_timer.N_382\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__41160\,
            I => \delay_measurement_inst.delay_tr_timer.N_382\
        );

    \I__8876\ : InMux
    port map (
            O => \N__41155\,
            I => \N__41152\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__41152\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16\
        );

    \I__8874\ : InMux
    port map (
            O => \N__41149\,
            I => \N__41146\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__41146\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\
        );

    \I__8872\ : CascadeMux
    port map (
            O => \N__41143\,
            I => \N__41140\
        );

    \I__8871\ : InMux
    port map (
            O => \N__41140\,
            I => \N__41135\
        );

    \I__8870\ : CascadeMux
    port map (
            O => \N__41139\,
            I => \N__41132\
        );

    \I__8869\ : InMux
    port map (
            O => \N__41138\,
            I => \N__41129\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__41135\,
            I => \N__41126\
        );

    \I__8867\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41122\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__41129\,
            I => \N__41117\
        );

    \I__8865\ : Span4Mux_h
    port map (
            O => \N__41126\,
            I => \N__41117\
        );

    \I__8864\ : InMux
    port map (
            O => \N__41125\,
            I => \N__41114\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__41122\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__8862\ : Odrv4
    port map (
            O => \N__41117\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__41114\,
            I => \elapsed_time_ns_1_RNIDH2591_0_5\
        );

    \I__8860\ : CascadeMux
    port map (
            O => \N__41107\,
            I => \elapsed_time_ns_1_RNIA965M1_0_18_cascade_\
        );

    \I__8859\ : CascadeMux
    port map (
            O => \N__41104\,
            I => \N__41101\
        );

    \I__8858\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41097\
        );

    \I__8857\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41093\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__41097\,
            I => \N__41090\
        );

    \I__8855\ : InMux
    port map (
            O => \N__41096\,
            I => \N__41086\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__41093\,
            I => \N__41083\
        );

    \I__8853\ : Span4Mux_v
    port map (
            O => \N__41090\,
            I => \N__41080\
        );

    \I__8852\ : InMux
    port map (
            O => \N__41089\,
            I => \N__41077\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__41086\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__8850\ : Odrv4
    port map (
            O => \N__41083\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__8849\ : Odrv4
    port map (
            O => \N__41080\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__41077\,
            I => \elapsed_time_ns_1_RNICG2591_0_4\
        );

    \I__8847\ : InMux
    port map (
            O => \N__41068\,
            I => \N__41065\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__41065\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2\
        );

    \I__8845\ : CascadeMux
    port map (
            O => \N__41062\,
            I => \N__41057\
        );

    \I__8844\ : CascadeMux
    port map (
            O => \N__41061\,
            I => \N__41051\
        );

    \I__8843\ : CascadeMux
    port map (
            O => \N__41060\,
            I => \N__41046\
        );

    \I__8842\ : InMux
    port map (
            O => \N__41057\,
            I => \N__41036\
        );

    \I__8841\ : InMux
    port map (
            O => \N__41056\,
            I => \N__41026\
        );

    \I__8840\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41019\
        );

    \I__8839\ : InMux
    port map (
            O => \N__41054\,
            I => \N__41014\
        );

    \I__8838\ : InMux
    port map (
            O => \N__41051\,
            I => \N__41014\
        );

    \I__8837\ : CascadeMux
    port map (
            O => \N__41050\,
            I => \N__41011\
        );

    \I__8836\ : CascadeMux
    port map (
            O => \N__41049\,
            I => \N__41008\
        );

    \I__8835\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41004\
        );

    \I__8834\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41001\
        );

    \I__8833\ : InMux
    port map (
            O => \N__41044\,
            I => \N__40998\
        );

    \I__8832\ : InMux
    port map (
            O => \N__41043\,
            I => \N__40987\
        );

    \I__8831\ : InMux
    port map (
            O => \N__41042\,
            I => \N__40987\
        );

    \I__8830\ : InMux
    port map (
            O => \N__41041\,
            I => \N__40987\
        );

    \I__8829\ : InMux
    port map (
            O => \N__41040\,
            I => \N__40987\
        );

    \I__8828\ : InMux
    port map (
            O => \N__41039\,
            I => \N__40987\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__41036\,
            I => \N__40984\
        );

    \I__8826\ : InMux
    port map (
            O => \N__41035\,
            I => \N__40975\
        );

    \I__8825\ : InMux
    port map (
            O => \N__41034\,
            I => \N__40975\
        );

    \I__8824\ : InMux
    port map (
            O => \N__41033\,
            I => \N__40975\
        );

    \I__8823\ : InMux
    port map (
            O => \N__41032\,
            I => \N__40975\
        );

    \I__8822\ : CascadeMux
    port map (
            O => \N__41031\,
            I => \N__40969\
        );

    \I__8821\ : CascadeMux
    port map (
            O => \N__41030\,
            I => \N__40966\
        );

    \I__8820\ : CascadeMux
    port map (
            O => \N__41029\,
            I => \N__40963\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__41026\,
            I => \N__40960\
        );

    \I__8818\ : InMux
    port map (
            O => \N__41025\,
            I => \N__40951\
        );

    \I__8817\ : InMux
    port map (
            O => \N__41024\,
            I => \N__40951\
        );

    \I__8816\ : InMux
    port map (
            O => \N__41023\,
            I => \N__40951\
        );

    \I__8815\ : InMux
    port map (
            O => \N__41022\,
            I => \N__40951\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__41019\,
            I => \N__40946\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__41014\,
            I => \N__40946\
        );

    \I__8812\ : InMux
    port map (
            O => \N__41011\,
            I => \N__40943\
        );

    \I__8811\ : InMux
    port map (
            O => \N__41008\,
            I => \N__40938\
        );

    \I__8810\ : InMux
    port map (
            O => \N__41007\,
            I => \N__40938\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__41004\,
            I => \N__40929\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__41001\,
            I => \N__40929\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__40998\,
            I => \N__40929\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__40987\,
            I => \N__40929\
        );

    \I__8805\ : Span4Mux_v
    port map (
            O => \N__40984\,
            I => \N__40924\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__40975\,
            I => \N__40924\
        );

    \I__8803\ : InMux
    port map (
            O => \N__40974\,
            I => \N__40917\
        );

    \I__8802\ : InMux
    port map (
            O => \N__40973\,
            I => \N__40917\
        );

    \I__8801\ : InMux
    port map (
            O => \N__40972\,
            I => \N__40917\
        );

    \I__8800\ : InMux
    port map (
            O => \N__40969\,
            I => \N__40910\
        );

    \I__8799\ : InMux
    port map (
            O => \N__40966\,
            I => \N__40910\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40963\,
            I => \N__40910\
        );

    \I__8797\ : Odrv4
    port map (
            O => \N__40960\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__40951\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__8795\ : Odrv4
    port map (
            O => \N__40946\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40943\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__40938\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__8792\ : Odrv4
    port map (
            O => \N__40929\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__8791\ : Odrv4
    port map (
            O => \N__40924\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__40917\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__40910\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\
        );

    \I__8788\ : CascadeMux
    port map (
            O => \N__40891\,
            I => \elapsed_time_ns_1_RNI9865M1_0_17_cascade_\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40885\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__40885\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40882\,
            I => \N__40879\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__40879\,
            I => \N__40876\
        );

    \I__8783\ : Span4Mux_v
    port map (
            O => \N__40876\,
            I => \N__40873\
        );

    \I__8782\ : Odrv4
    port map (
            O => \N__40873\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40870\,
            I => \N__40867\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__40867\,
            I => \N__40864\
        );

    \I__8779\ : Odrv4
    port map (
            O => \N__40864\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5\
        );

    \I__8778\ : InMux
    port map (
            O => \N__40861\,
            I => \N__40858\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__40858\,
            I => \N__40853\
        );

    \I__8776\ : InMux
    port map (
            O => \N__40857\,
            I => \N__40848\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40856\,
            I => \N__40848\
        );

    \I__8774\ : Odrv4
    port map (
            O => \N__40853\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lt31_0_2\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__40848\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lt31_0_2\
        );

    \I__8772\ : CascadeMux
    port map (
            O => \N__40843\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4_cascade_\
        );

    \I__8771\ : CascadeMux
    port map (
            O => \N__40840\,
            I => \N__40836\
        );

    \I__8770\ : InMux
    port map (
            O => \N__40839\,
            I => \N__40832\
        );

    \I__8769\ : InMux
    port map (
            O => \N__40836\,
            I => \N__40827\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40835\,
            I => \N__40827\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__40832\,
            I => \delay_measurement_inst.delay_tr_timer.N_358\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__40827\,
            I => \delay_measurement_inst.delay_tr_timer.N_358\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40822\,
            I => \N__40810\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40821\,
            I => \N__40810\
        );

    \I__8763\ : InMux
    port map (
            O => \N__40820\,
            I => \N__40807\
        );

    \I__8762\ : InMux
    port map (
            O => \N__40819\,
            I => \N__40804\
        );

    \I__8761\ : CascadeMux
    port map (
            O => \N__40818\,
            I => \N__40801\
        );

    \I__8760\ : CascadeMux
    port map (
            O => \N__40817\,
            I => \N__40798\
        );

    \I__8759\ : CascadeMux
    port map (
            O => \N__40816\,
            I => \N__40795\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__40815\,
            I => \N__40792\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__40810\,
            I => \N__40789\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__40807\,
            I => \N__40771\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__40804\,
            I => \N__40771\
        );

    \I__8754\ : InMux
    port map (
            O => \N__40801\,
            I => \N__40768\
        );

    \I__8753\ : InMux
    port map (
            O => \N__40798\,
            I => \N__40761\
        );

    \I__8752\ : InMux
    port map (
            O => \N__40795\,
            I => \N__40761\
        );

    \I__8751\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40761\
        );

    \I__8750\ : Span4Mux_v
    port map (
            O => \N__40789\,
            I => \N__40758\
        );

    \I__8749\ : InMux
    port map (
            O => \N__40788\,
            I => \N__40755\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40787\,
            I => \N__40750\
        );

    \I__8747\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40750\
        );

    \I__8746\ : InMux
    port map (
            O => \N__40785\,
            I => \N__40745\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40745\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40783\,
            I => \N__40740\
        );

    \I__8743\ : InMux
    port map (
            O => \N__40782\,
            I => \N__40740\
        );

    \I__8742\ : InMux
    port map (
            O => \N__40781\,
            I => \N__40733\
        );

    \I__8741\ : InMux
    port map (
            O => \N__40780\,
            I => \N__40733\
        );

    \I__8740\ : InMux
    port map (
            O => \N__40779\,
            I => \N__40733\
        );

    \I__8739\ : InMux
    port map (
            O => \N__40778\,
            I => \N__40726\
        );

    \I__8738\ : InMux
    port map (
            O => \N__40777\,
            I => \N__40726\
        );

    \I__8737\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40726\
        );

    \I__8736\ : Odrv4
    port map (
            O => \N__40771\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__40768\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__40761\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8733\ : Odrv4
    port map (
            O => \N__40758\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__40755\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__40750\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__40745\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__40740\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__40733\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__40726\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40705\,
            I => \N__40702\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__40702\,
            I => \delay_measurement_inst.delay_tr_timer.N_354\
        );

    \I__8724\ : CascadeMux
    port map (
            O => \N__40699\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\
        );

    \I__8723\ : InMux
    port map (
            O => \N__40696\,
            I => \N__40693\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__40693\,
            I => \N__40689\
        );

    \I__8721\ : InMux
    port map (
            O => \N__40692\,
            I => \N__40686\
        );

    \I__8720\ : Span4Mux_v
    port map (
            O => \N__40689\,
            I => \N__40681\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__40686\,
            I => \N__40678\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40685\,
            I => \N__40675\
        );

    \I__8717\ : InMux
    port map (
            O => \N__40684\,
            I => \N__40671\
        );

    \I__8716\ : Span4Mux_h
    port map (
            O => \N__40681\,
            I => \N__40668\
        );

    \I__8715\ : Span4Mux_v
    port map (
            O => \N__40678\,
            I => \N__40663\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__40675\,
            I => \N__40663\
        );

    \I__8713\ : InMux
    port map (
            O => \N__40674\,
            I => \N__40660\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__40671\,
            I => \elapsed_time_ns_1_RNIK8NQL1_0_3\
        );

    \I__8711\ : Odrv4
    port map (
            O => \N__40668\,
            I => \elapsed_time_ns_1_RNIK8NQL1_0_3\
        );

    \I__8710\ : Odrv4
    port map (
            O => \N__40663\,
            I => \elapsed_time_ns_1_RNIK8NQL1_0_3\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__40660\,
            I => \elapsed_time_ns_1_RNIK8NQL1_0_3\
        );

    \I__8708\ : InMux
    port map (
            O => \N__40651\,
            I => \N__40648\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__40648\,
            I => \N__40645\
        );

    \I__8706\ : Odrv4
    port map (
            O => \N__40645\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6\
        );

    \I__8705\ : CascadeMux
    port map (
            O => \N__40642\,
            I => \N__40639\
        );

    \I__8704\ : InMux
    port map (
            O => \N__40639\,
            I => \N__40635\
        );

    \I__8703\ : InMux
    port map (
            O => \N__40638\,
            I => \N__40631\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__40635\,
            I => \N__40627\
        );

    \I__8701\ : InMux
    port map (
            O => \N__40634\,
            I => \N__40624\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__40631\,
            I => \N__40621\
        );

    \I__8699\ : InMux
    port map (
            O => \N__40630\,
            I => \N__40618\
        );

    \I__8698\ : Span4Mux_v
    port map (
            O => \N__40627\,
            I => \N__40613\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__40624\,
            I => \N__40613\
        );

    \I__8696\ : Odrv4
    port map (
            O => \N__40621\,
            I => \elapsed_time_ns_1_RNINBNQL1_0_6\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__40618\,
            I => \elapsed_time_ns_1_RNINBNQL1_0_6\
        );

    \I__8694\ : Odrv4
    port map (
            O => \N__40613\,
            I => \elapsed_time_ns_1_RNINBNQL1_0_6\
        );

    \I__8693\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40603\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__40603\,
            I => \delay_measurement_inst.delay_tr_timer.N_353\
        );

    \I__8691\ : CascadeMux
    port map (
            O => \N__40600\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\
        );

    \I__8690\ : CascadeMux
    port map (
            O => \N__40597\,
            I => \N__40594\
        );

    \I__8689\ : InMux
    port map (
            O => \N__40594\,
            I => \N__40591\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__40591\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\
        );

    \I__8687\ : CascadeMux
    port map (
            O => \N__40588\,
            I => \N__40585\
        );

    \I__8686\ : InMux
    port map (
            O => \N__40585\,
            I => \N__40581\
        );

    \I__8685\ : InMux
    port map (
            O => \N__40584\,
            I => \N__40578\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__40581\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__40578\,
            I => \elapsed_time_ns_1_RNIUDIF91_0_24\
        );

    \I__8682\ : CascadeMux
    port map (
            O => \N__40573\,
            I => \delay_measurement_inst.delay_tr_timer.N_379_cascade_\
        );

    \I__8681\ : CascadeMux
    port map (
            O => \N__40570\,
            I => \delay_measurement_inst.delay_tr9_cascade_\
        );

    \I__8680\ : CascadeMux
    port map (
            O => \N__40567\,
            I => \N__40564\
        );

    \I__8679\ : InMux
    port map (
            O => \N__40564\,
            I => \N__40560\
        );

    \I__8678\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40557\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__40560\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__40557\,
            I => \elapsed_time_ns_1_RNIRBJF91_0_30\
        );

    \I__8675\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40545\
        );

    \I__8674\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40545\
        );

    \I__8673\ : InMux
    port map (
            O => \N__40550\,
            I => \N__40542\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__40545\,
            I => \N__40539\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__40542\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8670\ : Odrv12
    port map (
            O => \N__40539\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8669\ : InMux
    port map (
            O => \N__40534\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__8668\ : CascadeMux
    port map (
            O => \N__40531\,
            I => \N__40527\
        );

    \I__8667\ : CascadeMux
    port map (
            O => \N__40530\,
            I => \N__40524\
        );

    \I__8666\ : InMux
    port map (
            O => \N__40527\,
            I => \N__40518\
        );

    \I__8665\ : InMux
    port map (
            O => \N__40524\,
            I => \N__40518\
        );

    \I__8664\ : InMux
    port map (
            O => \N__40523\,
            I => \N__40515\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__40518\,
            I => \N__40512\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__40515\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8661\ : Odrv12
    port map (
            O => \N__40512\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8660\ : InMux
    port map (
            O => \N__40507\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__8659\ : CascadeMux
    port map (
            O => \N__40504\,
            I => \N__40501\
        );

    \I__8658\ : InMux
    port map (
            O => \N__40501\,
            I => \N__40497\
        );

    \I__8657\ : InMux
    port map (
            O => \N__40500\,
            I => \N__40494\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__40497\,
            I => \N__40491\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__40494\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8654\ : Odrv12
    port map (
            O => \N__40491\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8653\ : InMux
    port map (
            O => \N__40486\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__8652\ : InMux
    port map (
            O => \N__40483\,
            I => \N__40467\
        );

    \I__8651\ : InMux
    port map (
            O => \N__40482\,
            I => \N__40467\
        );

    \I__8650\ : InMux
    port map (
            O => \N__40481\,
            I => \N__40467\
        );

    \I__8649\ : InMux
    port map (
            O => \N__40480\,
            I => \N__40467\
        );

    \I__8648\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40444\
        );

    \I__8647\ : InMux
    port map (
            O => \N__40478\,
            I => \N__40444\
        );

    \I__8646\ : InMux
    port map (
            O => \N__40477\,
            I => \N__40444\
        );

    \I__8645\ : InMux
    port map (
            O => \N__40476\,
            I => \N__40444\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__40467\,
            I => \N__40437\
        );

    \I__8643\ : InMux
    port map (
            O => \N__40466\,
            I => \N__40432\
        );

    \I__8642\ : InMux
    port map (
            O => \N__40465\,
            I => \N__40432\
        );

    \I__8641\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40423\
        );

    \I__8640\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40423\
        );

    \I__8639\ : InMux
    port map (
            O => \N__40462\,
            I => \N__40423\
        );

    \I__8638\ : InMux
    port map (
            O => \N__40461\,
            I => \N__40423\
        );

    \I__8637\ : InMux
    port map (
            O => \N__40460\,
            I => \N__40414\
        );

    \I__8636\ : InMux
    port map (
            O => \N__40459\,
            I => \N__40414\
        );

    \I__8635\ : InMux
    port map (
            O => \N__40458\,
            I => \N__40414\
        );

    \I__8634\ : InMux
    port map (
            O => \N__40457\,
            I => \N__40414\
        );

    \I__8633\ : InMux
    port map (
            O => \N__40456\,
            I => \N__40405\
        );

    \I__8632\ : InMux
    port map (
            O => \N__40455\,
            I => \N__40405\
        );

    \I__8631\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40405\
        );

    \I__8630\ : InMux
    port map (
            O => \N__40453\,
            I => \N__40405\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__40444\,
            I => \N__40398\
        );

    \I__8628\ : InMux
    port map (
            O => \N__40443\,
            I => \N__40389\
        );

    \I__8627\ : InMux
    port map (
            O => \N__40442\,
            I => \N__40389\
        );

    \I__8626\ : InMux
    port map (
            O => \N__40441\,
            I => \N__40389\
        );

    \I__8625\ : InMux
    port map (
            O => \N__40440\,
            I => \N__40389\
        );

    \I__8624\ : Span4Mux_v
    port map (
            O => \N__40437\,
            I => \N__40382\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__40432\,
            I => \N__40382\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__40423\,
            I => \N__40382\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__40414\,
            I => \N__40379\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__40405\,
            I => \N__40376\
        );

    \I__8619\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40367\
        );

    \I__8618\ : InMux
    port map (
            O => \N__40403\,
            I => \N__40367\
        );

    \I__8617\ : InMux
    port map (
            O => \N__40402\,
            I => \N__40367\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40401\,
            I => \N__40367\
        );

    \I__8615\ : Span4Mux_v
    port map (
            O => \N__40398\,
            I => \N__40358\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__40389\,
            I => \N__40358\
        );

    \I__8613\ : Span4Mux_v
    port map (
            O => \N__40382\,
            I => \N__40358\
        );

    \I__8612\ : Span4Mux_v
    port map (
            O => \N__40379\,
            I => \N__40358\
        );

    \I__8611\ : Span4Mux_v
    port map (
            O => \N__40376\,
            I => \N__40353\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__40367\,
            I => \N__40353\
        );

    \I__8609\ : Span4Mux_h
    port map (
            O => \N__40358\,
            I => \N__40348\
        );

    \I__8608\ : Span4Mux_h
    port map (
            O => \N__40353\,
            I => \N__40348\
        );

    \I__8607\ : Odrv4
    port map (
            O => \N__40348\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8606\ : InMux
    port map (
            O => \N__40345\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__8605\ : InMux
    port map (
            O => \N__40342\,
            I => \N__40338\
        );

    \I__8604\ : InMux
    port map (
            O => \N__40341\,
            I => \N__40335\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__40338\,
            I => \N__40332\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__40335\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8601\ : Odrv12
    port map (
            O => \N__40332\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8600\ : CEMux
    port map (
            O => \N__40327\,
            I => \N__40322\
        );

    \I__8599\ : CEMux
    port map (
            O => \N__40326\,
            I => \N__40319\
        );

    \I__8598\ : CEMux
    port map (
            O => \N__40325\,
            I => \N__40315\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__40322\,
            I => \N__40310\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__40319\,
            I => \N__40310\
        );

    \I__8595\ : CEMux
    port map (
            O => \N__40318\,
            I => \N__40307\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__40315\,
            I => \N__40304\
        );

    \I__8593\ : Span4Mux_v
    port map (
            O => \N__40310\,
            I => \N__40301\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__40307\,
            I => \N__40298\
        );

    \I__8591\ : Span4Mux_v
    port map (
            O => \N__40304\,
            I => \N__40291\
        );

    \I__8590\ : Span4Mux_h
    port map (
            O => \N__40301\,
            I => \N__40291\
        );

    \I__8589\ : Span4Mux_h
    port map (
            O => \N__40298\,
            I => \N__40291\
        );

    \I__8588\ : Span4Mux_h
    port map (
            O => \N__40291\,
            I => \N__40288\
        );

    \I__8587\ : Odrv4
    port map (
            O => \N__40288\,
            I => \delay_measurement_inst.delay_hc_timer.N_398_i\
        );

    \I__8586\ : InMux
    port map (
            O => \N__40285\,
            I => \N__40282\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__40282\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20\
        );

    \I__8584\ : InMux
    port map (
            O => \N__40279\,
            I => \N__40275\
        );

    \I__8583\ : InMux
    port map (
            O => \N__40278\,
            I => \N__40272\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__40275\,
            I => \elapsed_time_ns_1_RNIRAIF91_0_21\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40272\,
            I => \elapsed_time_ns_1_RNIRAIF91_0_21\
        );

    \I__8580\ : CascadeMux
    port map (
            O => \N__40267\,
            I => \elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_\
        );

    \I__8579\ : InMux
    port map (
            O => \N__40264\,
            I => \N__40258\
        );

    \I__8578\ : InMux
    port map (
            O => \N__40263\,
            I => \N__40258\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__40258\,
            I => \elapsed_time_ns_1_RNI3JIF91_0_29\
        );

    \I__8576\ : InMux
    port map (
            O => \N__40255\,
            I => \N__40252\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__40252\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15\
        );

    \I__8574\ : InMux
    port map (
            O => \N__40249\,
            I => \N__40246\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__40246\,
            I => \elapsed_time_ns_1_RNITCIF91_0_23\
        );

    \I__8572\ : InMux
    port map (
            O => \N__40243\,
            I => \N__40240\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__40240\,
            I => \N__40235\
        );

    \I__8570\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40232\
        );

    \I__8569\ : InMux
    port map (
            O => \N__40238\,
            I => \N__40229\
        );

    \I__8568\ : Span4Mux_h
    port map (
            O => \N__40235\,
            I => \N__40226\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__40232\,
            I => \N__40223\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__40229\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8565\ : Odrv4
    port map (
            O => \N__40226\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8564\ : Odrv12
    port map (
            O => \N__40223\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8563\ : InMux
    port map (
            O => \N__40216\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__8562\ : CascadeMux
    port map (
            O => \N__40213\,
            I => \N__40210\
        );

    \I__8561\ : InMux
    port map (
            O => \N__40210\,
            I => \N__40206\
        );

    \I__8560\ : InMux
    port map (
            O => \N__40209\,
            I => \N__40203\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__40206\,
            I => \N__40197\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__40203\,
            I => \N__40197\
        );

    \I__8557\ : InMux
    port map (
            O => \N__40202\,
            I => \N__40194\
        );

    \I__8556\ : Span4Mux_h
    port map (
            O => \N__40197\,
            I => \N__40191\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__40194\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__8554\ : Odrv4
    port map (
            O => \N__40191\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__8553\ : InMux
    port map (
            O => \N__40186\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__8552\ : CascadeMux
    port map (
            O => \N__40183\,
            I => \N__40179\
        );

    \I__8551\ : CascadeMux
    port map (
            O => \N__40182\,
            I => \N__40176\
        );

    \I__8550\ : InMux
    port map (
            O => \N__40179\,
            I => \N__40170\
        );

    \I__8549\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40170\
        );

    \I__8548\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40167\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__40170\,
            I => \N__40164\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__40167\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8545\ : Odrv12
    port map (
            O => \N__40164\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8544\ : InMux
    port map (
            O => \N__40159\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__8543\ : InMux
    port map (
            O => \N__40156\,
            I => \N__40149\
        );

    \I__8542\ : InMux
    port map (
            O => \N__40155\,
            I => \N__40149\
        );

    \I__8541\ : InMux
    port map (
            O => \N__40154\,
            I => \N__40146\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__40149\,
            I => \N__40143\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__40146\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8538\ : Odrv12
    port map (
            O => \N__40143\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8537\ : InMux
    port map (
            O => \N__40138\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__8536\ : CascadeMux
    port map (
            O => \N__40135\,
            I => \N__40132\
        );

    \I__8535\ : InMux
    port map (
            O => \N__40132\,
            I => \N__40127\
        );

    \I__8534\ : InMux
    port map (
            O => \N__40131\,
            I => \N__40124\
        );

    \I__8533\ : InMux
    port map (
            O => \N__40130\,
            I => \N__40121\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__40127\,
            I => \N__40116\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__40124\,
            I => \N__40116\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__40121\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8529\ : Odrv12
    port map (
            O => \N__40116\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8528\ : InMux
    port map (
            O => \N__40111\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__8527\ : CascadeMux
    port map (
            O => \N__40108\,
            I => \N__40104\
        );

    \I__8526\ : CascadeMux
    port map (
            O => \N__40107\,
            I => \N__40101\
        );

    \I__8525\ : InMux
    port map (
            O => \N__40104\,
            I => \N__40096\
        );

    \I__8524\ : InMux
    port map (
            O => \N__40101\,
            I => \N__40096\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__40096\,
            I => \N__40092\
        );

    \I__8522\ : InMux
    port map (
            O => \N__40095\,
            I => \N__40089\
        );

    \I__8521\ : Span4Mux_v
    port map (
            O => \N__40092\,
            I => \N__40086\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__40089\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8519\ : Odrv4
    port map (
            O => \N__40086\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8518\ : InMux
    port map (
            O => \N__40081\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__8517\ : InMux
    port map (
            O => \N__40078\,
            I => \N__40071\
        );

    \I__8516\ : InMux
    port map (
            O => \N__40077\,
            I => \N__40071\
        );

    \I__8515\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40068\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__40071\,
            I => \N__40065\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__40068\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8512\ : Odrv12
    port map (
            O => \N__40065\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8511\ : InMux
    port map (
            O => \N__40060\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__8510\ : CascadeMux
    port map (
            O => \N__40057\,
            I => \N__40054\
        );

    \I__8509\ : InMux
    port map (
            O => \N__40054\,
            I => \N__40051\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__40051\,
            I => \N__40046\
        );

    \I__8507\ : InMux
    port map (
            O => \N__40050\,
            I => \N__40043\
        );

    \I__8506\ : InMux
    port map (
            O => \N__40049\,
            I => \N__40040\
        );

    \I__8505\ : Span4Mux_h
    port map (
            O => \N__40046\,
            I => \N__40037\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__40043\,
            I => \N__40034\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__40040\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8502\ : Odrv4
    port map (
            O => \N__40037\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8501\ : Odrv12
    port map (
            O => \N__40034\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8500\ : InMux
    port map (
            O => \N__40027\,
            I => \bfn_15_24_0_\
        );

    \I__8499\ : InMux
    port map (
            O => \N__40024\,
            I => \N__40020\
        );

    \I__8498\ : CascadeMux
    port map (
            O => \N__40023\,
            I => \N__40017\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__40020\,
            I => \N__40013\
        );

    \I__8496\ : InMux
    port map (
            O => \N__40017\,
            I => \N__40010\
        );

    \I__8495\ : InMux
    port map (
            O => \N__40016\,
            I => \N__40007\
        );

    \I__8494\ : Span4Mux_h
    port map (
            O => \N__40013\,
            I => \N__40004\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__40010\,
            I => \N__40001\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__40007\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8491\ : Odrv4
    port map (
            O => \N__40004\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8490\ : Odrv12
    port map (
            O => \N__40001\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39994\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__8488\ : CascadeMux
    port map (
            O => \N__39991\,
            I => \N__39988\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39988\,
            I => \N__39984\
        );

    \I__8486\ : InMux
    port map (
            O => \N__39987\,
            I => \N__39981\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__39984\,
            I => \N__39975\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__39981\,
            I => \N__39975\
        );

    \I__8483\ : InMux
    port map (
            O => \N__39980\,
            I => \N__39972\
        );

    \I__8482\ : Span4Mux_v
    port map (
            O => \N__39975\,
            I => \N__39969\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__39972\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__8480\ : Odrv4
    port map (
            O => \N__39969\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__8479\ : InMux
    port map (
            O => \N__39964\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__8478\ : InMux
    port map (
            O => \N__39961\,
            I => \N__39955\
        );

    \I__8477\ : InMux
    port map (
            O => \N__39960\,
            I => \N__39955\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39955\,
            I => \N__39951\
        );

    \I__8475\ : InMux
    port map (
            O => \N__39954\,
            I => \N__39948\
        );

    \I__8474\ : Span4Mux_h
    port map (
            O => \N__39951\,
            I => \N__39945\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__39948\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__8472\ : Odrv4
    port map (
            O => \N__39945\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39940\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39937\,
            I => \N__39931\
        );

    \I__8469\ : InMux
    port map (
            O => \N__39936\,
            I => \N__39931\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__39931\,
            I => \N__39927\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39924\
        );

    \I__8466\ : Span4Mux_h
    port map (
            O => \N__39927\,
            I => \N__39921\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__39924\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__8464\ : Odrv4
    port map (
            O => \N__39921\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__8463\ : InMux
    port map (
            O => \N__39916\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__8462\ : CascadeMux
    port map (
            O => \N__39913\,
            I => \N__39909\
        );

    \I__8461\ : CascadeMux
    port map (
            O => \N__39912\,
            I => \N__39906\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39909\,
            I => \N__39901\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39906\,
            I => \N__39901\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__39901\,
            I => \N__39897\
        );

    \I__8457\ : InMux
    port map (
            O => \N__39900\,
            I => \N__39894\
        );

    \I__8456\ : Span4Mux_v
    port map (
            O => \N__39897\,
            I => \N__39891\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__39894\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__39891\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__8453\ : InMux
    port map (
            O => \N__39886\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__8452\ : CascadeMux
    port map (
            O => \N__39883\,
            I => \N__39879\
        );

    \I__8451\ : CascadeMux
    port map (
            O => \N__39882\,
            I => \N__39876\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39879\,
            I => \N__39871\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39876\,
            I => \N__39871\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39871\,
            I => \N__39867\
        );

    \I__8447\ : InMux
    port map (
            O => \N__39870\,
            I => \N__39864\
        );

    \I__8446\ : Span4Mux_h
    port map (
            O => \N__39867\,
            I => \N__39861\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39864\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__8444\ : Odrv4
    port map (
            O => \N__39861\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39856\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__8442\ : CascadeMux
    port map (
            O => \N__39853\,
            I => \N__39850\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39850\,
            I => \N__39846\
        );

    \I__8440\ : InMux
    port map (
            O => \N__39849\,
            I => \N__39843\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__39846\,
            I => \N__39837\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__39843\,
            I => \N__39837\
        );

    \I__8437\ : InMux
    port map (
            O => \N__39842\,
            I => \N__39834\
        );

    \I__8436\ : Span4Mux_v
    port map (
            O => \N__39837\,
            I => \N__39831\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__39834\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__39831\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39826\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__8432\ : CascadeMux
    port map (
            O => \N__39823\,
            I => \N__39820\
        );

    \I__8431\ : InMux
    port map (
            O => \N__39820\,
            I => \N__39816\
        );

    \I__8430\ : InMux
    port map (
            O => \N__39819\,
            I => \N__39813\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__39816\,
            I => \N__39807\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__39813\,
            I => \N__39807\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39804\
        );

    \I__8426\ : Span4Mux_v
    port map (
            O => \N__39807\,
            I => \N__39801\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__39804\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__8424\ : Odrv4
    port map (
            O => \N__39801\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__8423\ : InMux
    port map (
            O => \N__39796\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__8422\ : CascadeMux
    port map (
            O => \N__39793\,
            I => \N__39790\
        );

    \I__8421\ : InMux
    port map (
            O => \N__39790\,
            I => \N__39786\
        );

    \I__8420\ : InMux
    port map (
            O => \N__39789\,
            I => \N__39783\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__39786\,
            I => \N__39779\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__39783\,
            I => \N__39776\
        );

    \I__8417\ : InMux
    port map (
            O => \N__39782\,
            I => \N__39773\
        );

    \I__8416\ : Span4Mux_v
    port map (
            O => \N__39779\,
            I => \N__39768\
        );

    \I__8415\ : Span4Mux_v
    port map (
            O => \N__39776\,
            I => \N__39768\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__39773\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__8413\ : Odrv4
    port map (
            O => \N__39768\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39763\,
            I => \bfn_15_23_0_\
        );

    \I__8411\ : CascadeMux
    port map (
            O => \N__39760\,
            I => \N__39756\
        );

    \I__8410\ : InMux
    port map (
            O => \N__39759\,
            I => \N__39753\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39756\,
            I => \N__39750\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__39753\,
            I => \N__39747\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__39750\,
            I => \N__39743\
        );

    \I__8406\ : Span4Mux_h
    port map (
            O => \N__39747\,
            I => \N__39740\
        );

    \I__8405\ : InMux
    port map (
            O => \N__39746\,
            I => \N__39737\
        );

    \I__8404\ : Span4Mux_h
    port map (
            O => \N__39743\,
            I => \N__39734\
        );

    \I__8403\ : Odrv4
    port map (
            O => \N__39740\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__39737\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8401\ : Odrv4
    port map (
            O => \N__39734\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8400\ : InMux
    port map (
            O => \N__39727\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__8399\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39717\
        );

    \I__8398\ : InMux
    port map (
            O => \N__39723\,
            I => \N__39717\
        );

    \I__8397\ : InMux
    port map (
            O => \N__39722\,
            I => \N__39714\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__39717\,
            I => \N__39711\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__39714\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__8394\ : Odrv12
    port map (
            O => \N__39711\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__8393\ : InMux
    port map (
            O => \N__39706\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__8392\ : InMux
    port map (
            O => \N__39703\,
            I => \N__39697\
        );

    \I__8391\ : InMux
    port map (
            O => \N__39702\,
            I => \N__39697\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__39697\,
            I => \N__39693\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39696\,
            I => \N__39690\
        );

    \I__8388\ : Span4Mux_v
    port map (
            O => \N__39693\,
            I => \N__39687\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__39690\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__8386\ : Odrv4
    port map (
            O => \N__39687\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__8385\ : InMux
    port map (
            O => \N__39682\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__8384\ : CascadeMux
    port map (
            O => \N__39679\,
            I => \N__39675\
        );

    \I__8383\ : InMux
    port map (
            O => \N__39678\,
            I => \N__39671\
        );

    \I__8382\ : InMux
    port map (
            O => \N__39675\,
            I => \N__39668\
        );

    \I__8381\ : InMux
    port map (
            O => \N__39674\,
            I => \N__39665\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__39671\,
            I => \N__39660\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__39668\,
            I => \N__39660\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__39665\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__8377\ : Odrv12
    port map (
            O => \N__39660\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__8376\ : InMux
    port map (
            O => \N__39655\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__8375\ : CascadeMux
    port map (
            O => \N__39652\,
            I => \N__39648\
        );

    \I__8374\ : CascadeMux
    port map (
            O => \N__39651\,
            I => \N__39645\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39648\,
            I => \N__39640\
        );

    \I__8372\ : InMux
    port map (
            O => \N__39645\,
            I => \N__39640\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__39640\,
            I => \N__39636\
        );

    \I__8370\ : InMux
    port map (
            O => \N__39639\,
            I => \N__39633\
        );

    \I__8369\ : Span4Mux_h
    port map (
            O => \N__39636\,
            I => \N__39630\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__39633\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__8367\ : Odrv4
    port map (
            O => \N__39630\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__8366\ : InMux
    port map (
            O => \N__39625\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__8365\ : CascadeMux
    port map (
            O => \N__39622\,
            I => \N__39618\
        );

    \I__8364\ : CascadeMux
    port map (
            O => \N__39621\,
            I => \N__39615\
        );

    \I__8363\ : InMux
    port map (
            O => \N__39618\,
            I => \N__39610\
        );

    \I__8362\ : InMux
    port map (
            O => \N__39615\,
            I => \N__39610\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__39610\,
            I => \N__39606\
        );

    \I__8360\ : InMux
    port map (
            O => \N__39609\,
            I => \N__39603\
        );

    \I__8359\ : Span4Mux_v
    port map (
            O => \N__39606\,
            I => \N__39600\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__39603\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__8357\ : Odrv4
    port map (
            O => \N__39600\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__8356\ : InMux
    port map (
            O => \N__39595\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__8355\ : CascadeMux
    port map (
            O => \N__39592\,
            I => \N__39589\
        );

    \I__8354\ : InMux
    port map (
            O => \N__39589\,
            I => \N__39585\
        );

    \I__8353\ : InMux
    port map (
            O => \N__39588\,
            I => \N__39582\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__39585\,
            I => \N__39576\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__39582\,
            I => \N__39576\
        );

    \I__8350\ : InMux
    port map (
            O => \N__39581\,
            I => \N__39573\
        );

    \I__8349\ : Span4Mux_v
    port map (
            O => \N__39576\,
            I => \N__39570\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__39573\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__8347\ : Odrv4
    port map (
            O => \N__39570\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__8346\ : InMux
    port map (
            O => \N__39565\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__39562\,
            I => \N__39559\
        );

    \I__8344\ : InMux
    port map (
            O => \N__39559\,
            I => \N__39556\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__39556\,
            I => \N__39551\
        );

    \I__8342\ : InMux
    port map (
            O => \N__39555\,
            I => \N__39548\
        );

    \I__8341\ : InMux
    port map (
            O => \N__39554\,
            I => \N__39545\
        );

    \I__8340\ : Span4Mux_h
    port map (
            O => \N__39551\,
            I => \N__39542\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__39548\,
            I => \N__39539\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__39545\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__8337\ : Odrv4
    port map (
            O => \N__39542\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__8336\ : Odrv12
    port map (
            O => \N__39539\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__8335\ : InMux
    port map (
            O => \N__39532\,
            I => \bfn_15_22_0_\
        );

    \I__8334\ : InMux
    port map (
            O => \N__39529\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__8333\ : InMux
    port map (
            O => \N__39526\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__8332\ : InMux
    port map (
            O => \N__39523\,
            I => \bfn_15_20_0_\
        );

    \I__8331\ : InMux
    port map (
            O => \N__39520\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__8330\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39513\
        );

    \I__8329\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39510\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__39513\,
            I => \N__39507\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__39510\,
            I => \N__39504\
        );

    \I__8326\ : Span4Mux_v
    port map (
            O => \N__39507\,
            I => \N__39499\
        );

    \I__8325\ : Span4Mux_h
    port map (
            O => \N__39504\,
            I => \N__39499\
        );

    \I__8324\ : Odrv4
    port map (
            O => \N__39499\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__8323\ : InMux
    port map (
            O => \N__39496\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__8322\ : CascadeMux
    port map (
            O => \N__39493\,
            I => \N__39490\
        );

    \I__8321\ : InMux
    port map (
            O => \N__39490\,
            I => \N__39486\
        );

    \I__8320\ : InMux
    port map (
            O => \N__39489\,
            I => \N__39483\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__39486\,
            I => \N__39480\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__39483\,
            I => \N__39477\
        );

    \I__8317\ : Span4Mux_h
    port map (
            O => \N__39480\,
            I => \N__39474\
        );

    \I__8316\ : Odrv12
    port map (
            O => \N__39477\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__8315\ : Odrv4
    port map (
            O => \N__39474\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__8314\ : InMux
    port map (
            O => \N__39469\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__8313\ : InMux
    port map (
            O => \N__39466\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__8312\ : InMux
    port map (
            O => \N__39463\,
            I => \N__39460\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__39460\,
            I => \N__39457\
        );

    \I__8310\ : Span4Mux_h
    port map (
            O => \N__39457\,
            I => \N__39454\
        );

    \I__8309\ : Odrv4
    port map (
            O => \N__39454\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__8308\ : CEMux
    port map (
            O => \N__39451\,
            I => \N__39436\
        );

    \I__8307\ : CEMux
    port map (
            O => \N__39450\,
            I => \N__39436\
        );

    \I__8306\ : CEMux
    port map (
            O => \N__39449\,
            I => \N__39436\
        );

    \I__8305\ : CEMux
    port map (
            O => \N__39448\,
            I => \N__39436\
        );

    \I__8304\ : CEMux
    port map (
            O => \N__39447\,
            I => \N__39436\
        );

    \I__8303\ : GlobalMux
    port map (
            O => \N__39436\,
            I => \N__39433\
        );

    \I__8302\ : gio2CtrlBuf
    port map (
            O => \N__39433\,
            I => \delay_measurement_inst.delay_hc_timer.N_397_i_g\
        );

    \I__8301\ : CascadeMux
    port map (
            O => \N__39430\,
            I => \N__39427\
        );

    \I__8300\ : InMux
    port map (
            O => \N__39427\,
            I => \N__39424\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__39424\,
            I => \N__39419\
        );

    \I__8298\ : InMux
    port map (
            O => \N__39423\,
            I => \N__39416\
        );

    \I__8297\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39413\
        );

    \I__8296\ : Span4Mux_h
    port map (
            O => \N__39419\,
            I => \N__39410\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__39416\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__39413\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8293\ : Odrv4
    port map (
            O => \N__39410\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8292\ : InMux
    port map (
            O => \N__39403\,
            I => \bfn_15_21_0_\
        );

    \I__8291\ : InMux
    port map (
            O => \N__39400\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__8290\ : InMux
    port map (
            O => \N__39397\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__8289\ : InMux
    port map (
            O => \N__39394\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__8288\ : InMux
    port map (
            O => \N__39391\,
            I => \bfn_15_19_0_\
        );

    \I__8287\ : InMux
    port map (
            O => \N__39388\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__8286\ : InMux
    port map (
            O => \N__39385\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8285\ : InMux
    port map (
            O => \N__39382\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8284\ : InMux
    port map (
            O => \N__39379\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8283\ : InMux
    port map (
            O => \N__39376\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8282\ : InMux
    port map (
            O => \N__39373\,
            I => \N__39367\
        );

    \I__8281\ : InMux
    port map (
            O => \N__39372\,
            I => \N__39367\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__39367\,
            I => \N__39364\
        );

    \I__8279\ : Odrv4
    port map (
            O => \N__39364\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__8278\ : InMux
    port map (
            O => \N__39361\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__8277\ : InMux
    port map (
            O => \N__39358\,
            I => \N__39352\
        );

    \I__8276\ : InMux
    port map (
            O => \N__39357\,
            I => \N__39352\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__39352\,
            I => \N__39349\
        );

    \I__8274\ : Odrv12
    port map (
            O => \N__39349\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__8273\ : InMux
    port map (
            O => \N__39346\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__8272\ : InMux
    port map (
            O => \N__39343\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__8271\ : InMux
    port map (
            O => \N__39340\,
            I => \N__39336\
        );

    \I__8270\ : InMux
    port map (
            O => \N__39339\,
            I => \N__39333\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__39336\,
            I => \N__39330\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__39333\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__8267\ : Odrv4
    port map (
            O => \N__39330\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__8266\ : InMux
    port map (
            O => \N__39325\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__8265\ : InMux
    port map (
            O => \N__39322\,
            I => \bfn_15_18_0_\
        );

    \I__8264\ : InMux
    port map (
            O => \N__39319\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__8263\ : InMux
    port map (
            O => \N__39316\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8262\ : InMux
    port map (
            O => \N__39313\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__8261\ : InMux
    port map (
            O => \N__39310\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__8260\ : InMux
    port map (
            O => \N__39307\,
            I => \N__39304\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__39304\,
            I => \N__39300\
        );

    \I__8258\ : InMux
    port map (
            O => \N__39303\,
            I => \N__39297\
        );

    \I__8257\ : Span4Mux_h
    port map (
            O => \N__39300\,
            I => \N__39293\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__39297\,
            I => \N__39290\
        );

    \I__8255\ : CascadeMux
    port map (
            O => \N__39296\,
            I => \N__39287\
        );

    \I__8254\ : Span4Mux_h
    port map (
            O => \N__39293\,
            I => \N__39284\
        );

    \I__8253\ : Span4Mux_v
    port map (
            O => \N__39290\,
            I => \N__39281\
        );

    \I__8252\ : InMux
    port map (
            O => \N__39287\,
            I => \N__39278\
        );

    \I__8251\ : Odrv4
    port map (
            O => \N__39284\,
            I => \elapsed_time_ns_1_RNILGKEE1_0_4\
        );

    \I__8250\ : Odrv4
    port map (
            O => \N__39281\,
            I => \elapsed_time_ns_1_RNILGKEE1_0_4\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__39278\,
            I => \elapsed_time_ns_1_RNILGKEE1_0_4\
        );

    \I__8248\ : CascadeMux
    port map (
            O => \N__39271\,
            I => \elapsed_time_ns_1_RNILGKEE1_0_4_cascade_\
        );

    \I__8247\ : InMux
    port map (
            O => \N__39268\,
            I => \N__39265\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__39265\,
            I => \N__39262\
        );

    \I__8245\ : Odrv4
    port map (
            O => \N__39262\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2\
        );

    \I__8244\ : InMux
    port map (
            O => \N__39259\,
            I => \N__39253\
        );

    \I__8243\ : InMux
    port map (
            O => \N__39258\,
            I => \N__39253\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__39253\,
            I => \elapsed_time_ns_1_RNI4GU8E1_0_21\
        );

    \I__8241\ : InMux
    port map (
            O => \N__39250\,
            I => \N__39244\
        );

    \I__8240\ : InMux
    port map (
            O => \N__39249\,
            I => \N__39244\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__39244\,
            I => \elapsed_time_ns_1_RNICOU8E1_0_29\
        );

    \I__8238\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39237\
        );

    \I__8237\ : InMux
    port map (
            O => \N__39240\,
            I => \N__39234\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__39237\,
            I => \N__39229\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__39234\,
            I => \N__39229\
        );

    \I__8234\ : Span4Mux_h
    port map (
            O => \N__39229\,
            I => \N__39226\
        );

    \I__8233\ : Odrv4
    port map (
            O => \N__39226\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__8232\ : InMux
    port map (
            O => \N__39223\,
            I => \N__39220\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__39220\,
            I => \N__39216\
        );

    \I__8230\ : InMux
    port map (
            O => \N__39219\,
            I => \N__39213\
        );

    \I__8229\ : Span4Mux_h
    port map (
            O => \N__39216\,
            I => \N__39210\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__39213\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__8227\ : Odrv4
    port map (
            O => \N__39210\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__8226\ : InMux
    port map (
            O => \N__39205\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__8225\ : InMux
    port map (
            O => \N__39202\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__8224\ : InMux
    port map (
            O => \N__39199\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__8223\ : InMux
    port map (
            O => \N__39196\,
            I => \N__39193\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__39193\,
            I => \N__39190\
        );

    \I__8221\ : Span4Mux_h
    port map (
            O => \N__39190\,
            I => \N__39187\
        );

    \I__8220\ : Odrv4
    port map (
            O => \N__39187\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df22\
        );

    \I__8219\ : InMux
    port map (
            O => \N__39184\,
            I => \N__39181\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__39181\,
            I => \N__39178\
        );

    \I__8217\ : Span4Mux_v
    port map (
            O => \N__39178\,
            I => \N__39175\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__39175\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df24\
        );

    \I__8215\ : InMux
    port map (
            O => \N__39172\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28\
        );

    \I__8214\ : InMux
    port map (
            O => \N__39169\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__8213\ : CascadeMux
    port map (
            O => \N__39166\,
            I => \N__39162\
        );

    \I__8212\ : InMux
    port map (
            O => \N__39165\,
            I => \N__39157\
        );

    \I__8211\ : InMux
    port map (
            O => \N__39162\,
            I => \N__39157\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__39157\,
            I => \elapsed_time_ns_1_RNI4HV8E1_0_30\
        );

    \I__8209\ : CascadeMux
    port map (
            O => \N__39154\,
            I => \N__39151\
        );

    \I__8208\ : InMux
    port map (
            O => \N__39151\,
            I => \N__39148\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__39148\,
            I => \N__39145\
        );

    \I__8206\ : Odrv12
    port map (
            O => \N__39145\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__8205\ : InMux
    port map (
            O => \N__39142\,
            I => \N__39139\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__39139\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__8203\ : InMux
    port map (
            O => \N__39136\,
            I => \N__39133\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__39133\,
            I => \N__39130\
        );

    \I__8201\ : Odrv12
    port map (
            O => \N__39130\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__8200\ : CascadeMux
    port map (
            O => \N__39127\,
            I => \N__39124\
        );

    \I__8199\ : InMux
    port map (
            O => \N__39124\,
            I => \N__39121\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__39121\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__8197\ : InMux
    port map (
            O => \N__39118\,
            I => \N__39115\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__39115\,
            I => \N__39112\
        );

    \I__8195\ : Odrv12
    port map (
            O => \N__39112\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__8194\ : CascadeMux
    port map (
            O => \N__39109\,
            I => \N__39106\
        );

    \I__8193\ : InMux
    port map (
            O => \N__39106\,
            I => \N__39103\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__39103\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__8191\ : InMux
    port map (
            O => \N__39100\,
            I => \N__39097\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__39097\,
            I => \N__39094\
        );

    \I__8189\ : Odrv12
    port map (
            O => \N__39094\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__8188\ : CascadeMux
    port map (
            O => \N__39091\,
            I => \N__39088\
        );

    \I__8187\ : InMux
    port map (
            O => \N__39088\,
            I => \N__39085\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__39085\,
            I => \N__39082\
        );

    \I__8185\ : Odrv4
    port map (
            O => \N__39082\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__8184\ : InMux
    port map (
            O => \N__39079\,
            I => \N__39076\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__39076\,
            I => \N__39073\
        );

    \I__8182\ : Odrv12
    port map (
            O => \N__39073\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__8181\ : CascadeMux
    port map (
            O => \N__39070\,
            I => \N__39067\
        );

    \I__8180\ : InMux
    port map (
            O => \N__39067\,
            I => \N__39064\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__39064\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__8178\ : InMux
    port map (
            O => \N__39061\,
            I => \N__39058\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__39058\,
            I => \N__39055\
        );

    \I__8176\ : Span4Mux_v
    port map (
            O => \N__39055\,
            I => \N__39052\
        );

    \I__8175\ : Odrv4
    port map (
            O => \N__39052\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__8174\ : CascadeMux
    port map (
            O => \N__39049\,
            I => \N__39046\
        );

    \I__8173\ : InMux
    port map (
            O => \N__39046\,
            I => \N__39043\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__39043\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__8171\ : InMux
    port map (
            O => \N__39040\,
            I => \N__39037\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__39037\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__8169\ : CascadeMux
    port map (
            O => \N__39034\,
            I => \N__39031\
        );

    \I__8168\ : InMux
    port map (
            O => \N__39031\,
            I => \N__39028\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__39028\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__8166\ : InMux
    port map (
            O => \N__39025\,
            I => \N__39022\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__39022\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__8164\ : CascadeMux
    port map (
            O => \N__39019\,
            I => \N__39016\
        );

    \I__8163\ : InMux
    port map (
            O => \N__39016\,
            I => \N__39013\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__39013\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__8161\ : InMux
    port map (
            O => \N__39010\,
            I => \N__39007\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__39007\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__8159\ : CascadeMux
    port map (
            O => \N__39004\,
            I => \N__39001\
        );

    \I__8158\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38998\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__38998\,
            I => \N__38995\
        );

    \I__8156\ : Odrv4
    port map (
            O => \N__38995\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__8155\ : InMux
    port map (
            O => \N__38992\,
            I => \N__38989\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38989\,
            I => \N__38986\
        );

    \I__8153\ : Span4Mux_v
    port map (
            O => \N__38986\,
            I => \N__38983\
        );

    \I__8152\ : Odrv4
    port map (
            O => \N__38983\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__8151\ : CascadeMux
    port map (
            O => \N__38980\,
            I => \N__38977\
        );

    \I__8150\ : InMux
    port map (
            O => \N__38977\,
            I => \N__38974\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__38974\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38971\,
            I => \N__38968\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__38968\,
            I => \N__38965\
        );

    \I__8146\ : Span4Mux_h
    port map (
            O => \N__38965\,
            I => \N__38962\
        );

    \I__8145\ : Odrv4
    port map (
            O => \N__38962\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__8144\ : CascadeMux
    port map (
            O => \N__38959\,
            I => \N__38956\
        );

    \I__8143\ : InMux
    port map (
            O => \N__38956\,
            I => \N__38953\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__38953\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38950\,
            I => \N__38947\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__38947\,
            I => \N__38944\
        );

    \I__8139\ : Odrv12
    port map (
            O => \N__38944\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__8138\ : CascadeMux
    port map (
            O => \N__38941\,
            I => \N__38938\
        );

    \I__8137\ : InMux
    port map (
            O => \N__38938\,
            I => \N__38935\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__38935\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__8135\ : InMux
    port map (
            O => \N__38932\,
            I => \N__38929\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__38929\,
            I => \N__38926\
        );

    \I__8133\ : Odrv12
    port map (
            O => \N__38926\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__8132\ : CascadeMux
    port map (
            O => \N__38923\,
            I => \N__38920\
        );

    \I__8131\ : InMux
    port map (
            O => \N__38920\,
            I => \N__38917\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__38917\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__8129\ : CascadeMux
    port map (
            O => \N__38914\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38911\,
            I => \N__38904\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38910\,
            I => \N__38904\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38909\,
            I => \N__38901\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__38904\,
            I => \elapsed_time_ns_1_RNII6NQL1_0_1\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38901\,
            I => \elapsed_time_ns_1_RNII6NQL1_0_1\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38896\,
            I => \N__38892\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38895\,
            I => \N__38889\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__38892\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__38889\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\
        );

    \I__8119\ : CascadeMux
    port map (
            O => \N__38884\,
            I => \elapsed_time_ns_1_RNII6NQL1_0_1_cascade_\
        );

    \I__8118\ : InMux
    port map (
            O => \N__38881\,
            I => \N__38878\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__38878\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38875\,
            I => \N__38871\
        );

    \I__8115\ : InMux
    port map (
            O => \N__38874\,
            I => \N__38868\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38871\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__38868\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\
        );

    \I__8112\ : CascadeMux
    port map (
            O => \N__38863\,
            I => \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\
        );

    \I__8111\ : CascadeMux
    port map (
            O => \N__38860\,
            I => \N__38857\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38857\,
            I => \N__38852\
        );

    \I__8109\ : CascadeMux
    port map (
            O => \N__38856\,
            I => \N__38846\
        );

    \I__8108\ : CascadeMux
    port map (
            O => \N__38855\,
            I => \N__38840\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__38852\,
            I => \N__38834\
        );

    \I__8106\ : InMux
    port map (
            O => \N__38851\,
            I => \N__38829\
        );

    \I__8105\ : InMux
    port map (
            O => \N__38850\,
            I => \N__38829\
        );

    \I__8104\ : InMux
    port map (
            O => \N__38849\,
            I => \N__38824\
        );

    \I__8103\ : InMux
    port map (
            O => \N__38846\,
            I => \N__38824\
        );

    \I__8102\ : InMux
    port map (
            O => \N__38845\,
            I => \N__38819\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38844\,
            I => \N__38819\
        );

    \I__8100\ : InMux
    port map (
            O => \N__38843\,
            I => \N__38808\
        );

    \I__8099\ : InMux
    port map (
            O => \N__38840\,
            I => \N__38808\
        );

    \I__8098\ : InMux
    port map (
            O => \N__38839\,
            I => \N__38808\
        );

    \I__8097\ : InMux
    port map (
            O => \N__38838\,
            I => \N__38808\
        );

    \I__8096\ : InMux
    port map (
            O => \N__38837\,
            I => \N__38808\
        );

    \I__8095\ : Span4Mux_h
    port map (
            O => \N__38834\,
            I => \N__38805\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__38829\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__38824\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__38819\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__38808\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__8090\ : Odrv4
    port map (
            O => \N__38805\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38794\,
            I => \N__38783\
        );

    \I__8088\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38783\
        );

    \I__8087\ : InMux
    port map (
            O => \N__38792\,
            I => \N__38783\
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__38791\,
            I => \N__38777\
        );

    \I__8085\ : CascadeMux
    port map (
            O => \N__38790\,
            I => \N__38773\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__38783\,
            I => \N__38765\
        );

    \I__8083\ : InMux
    port map (
            O => \N__38782\,
            I => \N__38760\
        );

    \I__8082\ : InMux
    port map (
            O => \N__38781\,
            I => \N__38760\
        );

    \I__8081\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38757\
        );

    \I__8080\ : InMux
    port map (
            O => \N__38777\,
            I => \N__38752\
        );

    \I__8079\ : InMux
    port map (
            O => \N__38776\,
            I => \N__38752\
        );

    \I__8078\ : InMux
    port map (
            O => \N__38773\,
            I => \N__38747\
        );

    \I__8077\ : InMux
    port map (
            O => \N__38772\,
            I => \N__38747\
        );

    \I__8076\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38738\
        );

    \I__8075\ : InMux
    port map (
            O => \N__38770\,
            I => \N__38738\
        );

    \I__8074\ : InMux
    port map (
            O => \N__38769\,
            I => \N__38738\
        );

    \I__8073\ : InMux
    port map (
            O => \N__38768\,
            I => \N__38738\
        );

    \I__8072\ : Span4Mux_h
    port map (
            O => \N__38765\,
            I => \N__38735\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__38760\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__38757\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__38752\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__38747\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__38738\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__8066\ : Odrv4
    port map (
            O => \N__38735\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__38722\,
            I => \N__38719\
        );

    \I__8064\ : InMux
    port map (
            O => \N__38719\,
            I => \N__38716\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__38716\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__8062\ : InMux
    port map (
            O => \N__38713\,
            I => \N__38710\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__38710\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__38707\,
            I => \N__38704\
        );

    \I__8059\ : InMux
    port map (
            O => \N__38704\,
            I => \N__38701\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__38701\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__8057\ : InMux
    port map (
            O => \N__38698\,
            I => \N__38695\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__38695\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__8055\ : InMux
    port map (
            O => \N__38692\,
            I => \N__38689\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__38689\,
            I => \N__38685\
        );

    \I__8053\ : InMux
    port map (
            O => \N__38688\,
            I => \N__38680\
        );

    \I__8052\ : Span4Mux_v
    port map (
            O => \N__38685\,
            I => \N__38677\
        );

    \I__8051\ : InMux
    port map (
            O => \N__38684\,
            I => \N__38674\
        );

    \I__8050\ : InMux
    port map (
            O => \N__38683\,
            I => \N__38671\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__38680\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\
        );

    \I__8048\ : Odrv4
    port map (
            O => \N__38677\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__38674\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__38671\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__38662\,
            I => \delay_measurement_inst.delay_tr_timer.N_386_cascade_\
        );

    \I__8044\ : InMux
    port map (
            O => \N__38659\,
            I => \N__38656\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__38656\,
            I => \N__38652\
        );

    \I__8042\ : InMux
    port map (
            O => \N__38655\,
            I => \N__38649\
        );

    \I__8041\ : Odrv4
    port map (
            O => \N__38652\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__38649\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__38644\,
            I => \N__38640\
        );

    \I__8038\ : CascadeMux
    port map (
            O => \N__38643\,
            I => \N__38637\
        );

    \I__8037\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38634\
        );

    \I__8036\ : InMux
    port map (
            O => \N__38637\,
            I => \N__38631\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__38634\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__38631\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2\
        );

    \I__8033\ : CascadeMux
    port map (
            O => \N__38626\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2_cascade_\
        );

    \I__8032\ : InMux
    port map (
            O => \N__38623\,
            I => \N__38616\
        );

    \I__8031\ : InMux
    port map (
            O => \N__38622\,
            I => \N__38616\
        );

    \I__8030\ : InMux
    port map (
            O => \N__38621\,
            I => \N__38613\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__38616\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__38613\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\
        );

    \I__8027\ : InMux
    port map (
            O => \N__38608\,
            I => \N__38603\
        );

    \I__8026\ : InMux
    port map (
            O => \N__38607\,
            I => \N__38598\
        );

    \I__8025\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38598\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__38603\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__38598\,
            I => \elapsed_time_ns_1_RNIAE2591_0_2\
        );

    \I__8022\ : InMux
    port map (
            O => \N__38593\,
            I => \N__38590\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__38590\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1\
        );

    \I__8020\ : CascadeMux
    port map (
            O => \N__38587\,
            I => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\
        );

    \I__8019\ : InMux
    port map (
            O => \N__38584\,
            I => \N__38580\
        );

    \I__8018\ : InMux
    port map (
            O => \N__38583\,
            I => \N__38577\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__38580\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__38577\,
            I => \elapsed_time_ns_1_RNI0GIF91_0_26\
        );

    \I__8015\ : CascadeMux
    port map (
            O => \N__38572\,
            I => \N__38568\
        );

    \I__8014\ : CascadeMux
    port map (
            O => \N__38571\,
            I => \N__38565\
        );

    \I__8013\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38561\
        );

    \I__8012\ : InMux
    port map (
            O => \N__38565\,
            I => \N__38558\
        );

    \I__8011\ : InMux
    port map (
            O => \N__38564\,
            I => \N__38555\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__38561\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__38558\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__38555\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10\
        );

    \I__8007\ : InMux
    port map (
            O => \N__38548\,
            I => \N__38542\
        );

    \I__8006\ : InMux
    port map (
            O => \N__38547\,
            I => \N__38539\
        );

    \I__8005\ : InMux
    port map (
            O => \N__38546\,
            I => \N__38536\
        );

    \I__8004\ : InMux
    port map (
            O => \N__38545\,
            I => \N__38533\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__38542\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__38539\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__38536\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__38533\,
            I => \elapsed_time_ns_1_RNIQ8HF91_0_11\
        );

    \I__7999\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38518\
        );

    \I__7998\ : InMux
    port map (
            O => \N__38523\,
            I => \N__38515\
        );

    \I__7997\ : InMux
    port map (
            O => \N__38522\,
            I => \N__38512\
        );

    \I__7996\ : InMux
    port map (
            O => \N__38521\,
            I => \N__38509\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__38518\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__38515\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__38512\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__38509\,
            I => \elapsed_time_ns_1_RNIR9HF91_0_12\
        );

    \I__7991\ : CascadeMux
    port map (
            O => \N__38500\,
            I => \N__38496\
        );

    \I__7990\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38491\
        );

    \I__7989\ : InMux
    port map (
            O => \N__38496\,
            I => \N__38488\
        );

    \I__7988\ : InMux
    port map (
            O => \N__38495\,
            I => \N__38485\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38494\,
            I => \N__38482\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__38491\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__38488\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__38485\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__38482\,
            I => \elapsed_time_ns_1_RNISAHF91_0_13\
        );

    \I__7982\ : InMux
    port map (
            O => \N__38473\,
            I => \N__38462\
        );

    \I__7981\ : InMux
    port map (
            O => \N__38472\,
            I => \N__38462\
        );

    \I__7980\ : InMux
    port map (
            O => \N__38471\,
            I => \N__38459\
        );

    \I__7979\ : InMux
    port map (
            O => \N__38470\,
            I => \N__38456\
        );

    \I__7978\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38453\
        );

    \I__7977\ : InMux
    port map (
            O => \N__38468\,
            I => \N__38448\
        );

    \I__7976\ : InMux
    port map (
            O => \N__38467\,
            I => \N__38448\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__38462\,
            I => \N__38445\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__38459\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__38456\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__38453\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__38448\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7970\ : Odrv4
    port map (
            O => \N__38445\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15\
        );

    \I__7969\ : CascadeMux
    port map (
            O => \N__38434\,
            I => \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\
        );

    \I__7968\ : CascadeMux
    port map (
            O => \N__38431\,
            I => \N__38423\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__38430\,
            I => \N__38420\
        );

    \I__7966\ : InMux
    port map (
            O => \N__38429\,
            I => \N__38411\
        );

    \I__7965\ : InMux
    port map (
            O => \N__38428\,
            I => \N__38400\
        );

    \I__7964\ : InMux
    port map (
            O => \N__38427\,
            I => \N__38400\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38426\,
            I => \N__38400\
        );

    \I__7962\ : InMux
    port map (
            O => \N__38423\,
            I => \N__38400\
        );

    \I__7961\ : InMux
    port map (
            O => \N__38420\,
            I => \N__38400\
        );

    \I__7960\ : InMux
    port map (
            O => \N__38419\,
            I => \N__38387\
        );

    \I__7959\ : InMux
    port map (
            O => \N__38418\,
            I => \N__38387\
        );

    \I__7958\ : InMux
    port map (
            O => \N__38417\,
            I => \N__38387\
        );

    \I__7957\ : InMux
    port map (
            O => \N__38416\,
            I => \N__38387\
        );

    \I__7956\ : InMux
    port map (
            O => \N__38415\,
            I => \N__38387\
        );

    \I__7955\ : InMux
    port map (
            O => \N__38414\,
            I => \N__38387\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__38411\,
            I => \phase_controller_inst1.stoper_tr.N_244\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__38400\,
            I => \phase_controller_inst1.stoper_tr.N_244\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__38387\,
            I => \phase_controller_inst1.stoper_tr.N_244\
        );

    \I__7951\ : InMux
    port map (
            O => \N__38380\,
            I => \N__38377\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__38377\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\
        );

    \I__7949\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38371\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__38371\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25\
        );

    \I__7947\ : CascadeMux
    port map (
            O => \N__38368\,
            I => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\
        );

    \I__7946\ : InMux
    port map (
            O => \N__38365\,
            I => \N__38359\
        );

    \I__7945\ : InMux
    port map (
            O => \N__38364\,
            I => \N__38359\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__38359\,
            I => \elapsed_time_ns_1_RNI2IIF91_0_28\
        );

    \I__7943\ : CascadeMux
    port map (
            O => \N__38356\,
            I => \N__38353\
        );

    \I__7942\ : InMux
    port map (
            O => \N__38353\,
            I => \N__38347\
        );

    \I__7941\ : InMux
    port map (
            O => \N__38352\,
            I => \N__38347\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__38347\,
            I => \elapsed_time_ns_1_RNI1HIF91_0_27\
        );

    \I__7939\ : InMux
    port map (
            O => \N__38344\,
            I => \N__38341\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__38341\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15\
        );

    \I__7937\ : CascadeMux
    port map (
            O => \N__38338\,
            I => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_\
        );

    \I__7936\ : CascadeMux
    port map (
            O => \N__38335\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\
        );

    \I__7935\ : InMux
    port map (
            O => \N__38332\,
            I => \N__38326\
        );

    \I__7934\ : InMux
    port map (
            O => \N__38331\,
            I => \N__38326\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__38326\,
            I => \elapsed_time_ns_1_RNISBIF91_0_22\
        );

    \I__7932\ : CascadeMux
    port map (
            O => \N__38323\,
            I => \N__38319\
        );

    \I__7931\ : InMux
    port map (
            O => \N__38322\,
            I => \N__38316\
        );

    \I__7930\ : InMux
    port map (
            O => \N__38319\,
            I => \N__38313\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__38316\,
            I => \N__38309\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__38313\,
            I => \N__38306\
        );

    \I__7927\ : InMux
    port map (
            O => \N__38312\,
            I => \N__38303\
        );

    \I__7926\ : Odrv4
    port map (
            O => \N__38309\,
            I => \elapsed_time_ns_1_RNIOJKEE1_0_7\
        );

    \I__7925\ : Odrv4
    port map (
            O => \N__38306\,
            I => \elapsed_time_ns_1_RNIOJKEE1_0_7\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__38303\,
            I => \elapsed_time_ns_1_RNIOJKEE1_0_7\
        );

    \I__7923\ : CascadeMux
    port map (
            O => \N__38296\,
            I => \N__38291\
        );

    \I__7922\ : InMux
    port map (
            O => \N__38295\,
            I => \N__38288\
        );

    \I__7921\ : InMux
    port map (
            O => \N__38294\,
            I => \N__38285\
        );

    \I__7920\ : InMux
    port map (
            O => \N__38291\,
            I => \N__38282\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__38288\,
            I => \N__38279\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__38285\,
            I => \N__38274\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__38282\,
            I => \N__38274\
        );

    \I__7916\ : Span4Mux_h
    port map (
            O => \N__38279\,
            I => \N__38271\
        );

    \I__7915\ : Span12Mux_h
    port map (
            O => \N__38274\,
            I => \N__38266\
        );

    \I__7914\ : Sp12to4
    port map (
            O => \N__38271\,
            I => \N__38266\
        );

    \I__7913\ : Span12Mux_v
    port map (
            O => \N__38266\,
            I => \N__38263\
        );

    \I__7912\ : Odrv12
    port map (
            O => \N__38263\,
            I => \il_max_comp1_D2\
        );

    \I__7911\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38247\
        );

    \I__7910\ : InMux
    port map (
            O => \N__38259\,
            I => \N__38247\
        );

    \I__7909\ : InMux
    port map (
            O => \N__38258\,
            I => \N__38247\
        );

    \I__7908\ : InMux
    port map (
            O => \N__38257\,
            I => \N__38243\
        );

    \I__7907\ : InMux
    port map (
            O => \N__38256\,
            I => \N__38240\
        );

    \I__7906\ : InMux
    port map (
            O => \N__38255\,
            I => \N__38237\
        );

    \I__7905\ : InMux
    port map (
            O => \N__38254\,
            I => \N__38234\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__38247\,
            I => \N__38231\
        );

    \I__7903\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38228\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__38243\,
            I => state_3
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__38240\,
            I => state_3
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__38237\,
            I => state_3
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__38234\,
            I => state_3
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__38231\,
            I => state_3
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__38228\,
            I => state_3
        );

    \I__7896\ : IoInMux
    port map (
            O => \N__38215\,
            I => \N__38212\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__38212\,
            I => \N__38209\
        );

    \I__7894\ : IoSpan4Mux
    port map (
            O => \N__38209\,
            I => \N__38206\
        );

    \I__7893\ : Span4Mux_s3_v
    port map (
            O => \N__38206\,
            I => \N__38203\
        );

    \I__7892\ : Span4Mux_v
    port map (
            O => \N__38203\,
            I => \N__38199\
        );

    \I__7891\ : InMux
    port map (
            O => \N__38202\,
            I => \N__38196\
        );

    \I__7890\ : Odrv4
    port map (
            O => \N__38199\,
            I => \T01_c\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__38196\,
            I => \T01_c\
        );

    \I__7888\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38188\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__38188\,
            I => \N__38185\
        );

    \I__7886\ : Span4Mux_h
    port map (
            O => \N__38185\,
            I => \N__38182\
        );

    \I__7885\ : Odrv4
    port map (
            O => \N__38182\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__38179\,
            I => \N__38175\
        );

    \I__7883\ : CascadeMux
    port map (
            O => \N__38178\,
            I => \N__38171\
        );

    \I__7882\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38168\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__38174\,
            I => \N__38165\
        );

    \I__7880\ : InMux
    port map (
            O => \N__38171\,
            I => \N__38162\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__38168\,
            I => \N__38159\
        );

    \I__7878\ : InMux
    port map (
            O => \N__38165\,
            I => \N__38156\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__38162\,
            I => \N__38151\
        );

    \I__7876\ : Span4Mux_v
    port map (
            O => \N__38159\,
            I => \N__38146\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__38156\,
            I => \N__38146\
        );

    \I__7874\ : InMux
    port map (
            O => \N__38155\,
            I => \N__38141\
        );

    \I__7873\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38141\
        );

    \I__7872\ : Span4Mux_h
    port map (
            O => \N__38151\,
            I => \N__38138\
        );

    \I__7871\ : Span4Mux_h
    port map (
            O => \N__38146\,
            I => \N__38133\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__38141\,
            I => \N__38133\
        );

    \I__7869\ : Span4Mux_h
    port map (
            O => \N__38138\,
            I => \N__38130\
        );

    \I__7868\ : Span4Mux_h
    port map (
            O => \N__38133\,
            I => \N__38127\
        );

    \I__7867\ : Odrv4
    port map (
            O => \N__38130\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__7866\ : Odrv4
    port map (
            O => \N__38127\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__7865\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38119\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__38119\,
            I => \N__38116\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__38116\,
            I => \N__38113\
        );

    \I__7862\ : Odrv4
    port map (
            O => \N__38113\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__7861\ : CascadeMux
    port map (
            O => \N__38110\,
            I => \N__38107\
        );

    \I__7860\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38104\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__38104\,
            I => \N__38100\
        );

    \I__7858\ : InMux
    port map (
            O => \N__38103\,
            I => \N__38097\
        );

    \I__7857\ : Span4Mux_h
    port map (
            O => \N__38100\,
            I => \N__38090\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__38097\,
            I => \N__38090\
        );

    \I__7855\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38087\
        );

    \I__7854\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38083\
        );

    \I__7853\ : Span4Mux_v
    port map (
            O => \N__38090\,
            I => \N__38080\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__38087\,
            I => \N__38077\
        );

    \I__7851\ : InMux
    port map (
            O => \N__38086\,
            I => \N__38074\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__38083\,
            I => \N__38069\
        );

    \I__7849\ : Sp12to4
    port map (
            O => \N__38080\,
            I => \N__38069\
        );

    \I__7848\ : Span4Mux_h
    port map (
            O => \N__38077\,
            I => \N__38064\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__38074\,
            I => \N__38064\
        );

    \I__7846\ : Odrv12
    port map (
            O => \N__38069\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__7845\ : Odrv4
    port map (
            O => \N__38064\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__7844\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38054\
        );

    \I__7843\ : InMux
    port map (
            O => \N__38058\,
            I => \N__38051\
        );

    \I__7842\ : InMux
    port map (
            O => \N__38057\,
            I => \N__38048\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__38054\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__38051\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__38048\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\
        );

    \I__7838\ : CascadeMux
    port map (
            O => \N__38041\,
            I => \N__38038\
        );

    \I__7837\ : InMux
    port map (
            O => \N__38038\,
            I => \N__38032\
        );

    \I__7836\ : InMux
    port map (
            O => \N__38037\,
            I => \N__38029\
        );

    \I__7835\ : InMux
    port map (
            O => \N__38036\,
            I => \N__38026\
        );

    \I__7834\ : InMux
    port map (
            O => \N__38035\,
            I => \N__38023\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__38032\,
            I => \N__38020\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__38029\,
            I => \N__38017\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__38026\,
            I => \N__38014\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__38023\,
            I => \N__38011\
        );

    \I__7829\ : Span4Mux_v
    port map (
            O => \N__38020\,
            I => \N__38008\
        );

    \I__7828\ : Span4Mux_v
    port map (
            O => \N__38017\,
            I => \N__38005\
        );

    \I__7827\ : Span4Mux_h
    port map (
            O => \N__38014\,
            I => \N__38001\
        );

    \I__7826\ : Span4Mux_v
    port map (
            O => \N__38011\,
            I => \N__37994\
        );

    \I__7825\ : Span4Mux_h
    port map (
            O => \N__38008\,
            I => \N__37994\
        );

    \I__7824\ : Span4Mux_h
    port map (
            O => \N__38005\,
            I => \N__37994\
        );

    \I__7823\ : InMux
    port map (
            O => \N__38004\,
            I => \N__37991\
        );

    \I__7822\ : Odrv4
    port map (
            O => \N__38001\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__7821\ : Odrv4
    port map (
            O => \N__37994\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__37991\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__7819\ : CascadeMux
    port map (
            O => \N__37984\,
            I => \N__37980\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37983\,
            I => \N__37966\
        );

    \I__7817\ : InMux
    port map (
            O => \N__37980\,
            I => \N__37963\
        );

    \I__7816\ : InMux
    port map (
            O => \N__37979\,
            I => \N__37954\
        );

    \I__7815\ : InMux
    port map (
            O => \N__37978\,
            I => \N__37954\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37977\,
            I => \N__37954\
        );

    \I__7813\ : InMux
    port map (
            O => \N__37976\,
            I => \N__37954\
        );

    \I__7812\ : CascadeMux
    port map (
            O => \N__37975\,
            I => \N__37951\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37974\,
            I => \N__37919\
        );

    \I__7810\ : InMux
    port map (
            O => \N__37973\,
            I => \N__37919\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37972\,
            I => \N__37919\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37971\,
            I => \N__37919\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37970\,
            I => \N__37919\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37969\,
            I => \N__37919\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__37966\,
            I => \N__37916\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__37963\,
            I => \N__37911\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__37954\,
            I => \N__37911\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37951\,
            I => \N__37900\
        );

    \I__7801\ : InMux
    port map (
            O => \N__37950\,
            I => \N__37900\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37949\,
            I => \N__37900\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37900\
        );

    \I__7798\ : InMux
    port map (
            O => \N__37947\,
            I => \N__37900\
        );

    \I__7797\ : InMux
    port map (
            O => \N__37946\,
            I => \N__37897\
        );

    \I__7796\ : CascadeMux
    port map (
            O => \N__37945\,
            I => \N__37894\
        );

    \I__7795\ : CascadeMux
    port map (
            O => \N__37944\,
            I => \N__37889\
        );

    \I__7794\ : CascadeMux
    port map (
            O => \N__37943\,
            I => \N__37885\
        );

    \I__7793\ : CascadeMux
    port map (
            O => \N__37942\,
            I => \N__37879\
        );

    \I__7792\ : CascadeMux
    port map (
            O => \N__37941\,
            I => \N__37874\
        );

    \I__7791\ : CascadeMux
    port map (
            O => \N__37940\,
            I => \N__37868\
        );

    \I__7790\ : InMux
    port map (
            O => \N__37939\,
            I => \N__37860\
        );

    \I__7789\ : InMux
    port map (
            O => \N__37938\,
            I => \N__37860\
        );

    \I__7788\ : InMux
    port map (
            O => \N__37937\,
            I => \N__37860\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37936\,
            I => \N__37851\
        );

    \I__7786\ : InMux
    port map (
            O => \N__37935\,
            I => \N__37851\
        );

    \I__7785\ : InMux
    port map (
            O => \N__37934\,
            I => \N__37851\
        );

    \I__7784\ : InMux
    port map (
            O => \N__37933\,
            I => \N__37851\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37932\,
            I => \N__37848\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__37919\,
            I => \N__37839\
        );

    \I__7781\ : Span4Mux_v
    port map (
            O => \N__37916\,
            I => \N__37839\
        );

    \I__7780\ : Span4Mux_v
    port map (
            O => \N__37911\,
            I => \N__37839\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37900\,
            I => \N__37839\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__37897\,
            I => \N__37834\
        );

    \I__7777\ : InMux
    port map (
            O => \N__37894\,
            I => \N__37828\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37893\,
            I => \N__37828\
        );

    \I__7775\ : InMux
    port map (
            O => \N__37892\,
            I => \N__37817\
        );

    \I__7774\ : InMux
    port map (
            O => \N__37889\,
            I => \N__37817\
        );

    \I__7773\ : InMux
    port map (
            O => \N__37888\,
            I => \N__37817\
        );

    \I__7772\ : InMux
    port map (
            O => \N__37885\,
            I => \N__37817\
        );

    \I__7771\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37817\
        );

    \I__7770\ : InMux
    port map (
            O => \N__37883\,
            I => \N__37806\
        );

    \I__7769\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37806\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37879\,
            I => \N__37806\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37806\
        );

    \I__7766\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37806\
        );

    \I__7765\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37793\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37793\
        );

    \I__7763\ : InMux
    port map (
            O => \N__37872\,
            I => \N__37793\
        );

    \I__7762\ : InMux
    port map (
            O => \N__37871\,
            I => \N__37793\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37868\,
            I => \N__37793\
        );

    \I__7760\ : InMux
    port map (
            O => \N__37867\,
            I => \N__37793\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__37860\,
            I => \N__37786\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__37851\,
            I => \N__37786\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__37848\,
            I => \N__37781\
        );

    \I__7756\ : Span4Mux_h
    port map (
            O => \N__37839\,
            I => \N__37781\
        );

    \I__7755\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37776\
        );

    \I__7754\ : InMux
    port map (
            O => \N__37837\,
            I => \N__37776\
        );

    \I__7753\ : Span4Mux_h
    port map (
            O => \N__37834\,
            I => \N__37773\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37770\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__37828\,
            I => \N__37761\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__37817\,
            I => \N__37761\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__37806\,
            I => \N__37761\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__37793\,
            I => \N__37761\
        );

    \I__7747\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37756\
        );

    \I__7746\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37756\
        );

    \I__7745\ : Span4Mux_v
    port map (
            O => \N__37786\,
            I => \N__37751\
        );

    \I__7744\ : Span4Mux_v
    port map (
            O => \N__37781\,
            I => \N__37751\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__37776\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7742\ : Odrv4
    port map (
            O => \N__37773\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__37770\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7740\ : Odrv12
    port map (
            O => \N__37761\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__37756\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__37751\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7737\ : InMux
    port map (
            O => \N__37738\,
            I => \N__37735\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__37735\,
            I => \N__37732\
        );

    \I__7735\ : Odrv4
    port map (
            O => \N__37732\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\
        );

    \I__7734\ : CascadeMux
    port map (
            O => \N__37729\,
            I => \N__37726\
        );

    \I__7733\ : InMux
    port map (
            O => \N__37726\,
            I => \N__37723\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__37723\,
            I => \N__37720\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__37720\,
            I => \N__37717\
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__37717\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0\
        );

    \I__7729\ : CascadeMux
    port map (
            O => \N__37714\,
            I => \N__37710\
        );

    \I__7728\ : InMux
    port map (
            O => \N__37713\,
            I => \N__37703\
        );

    \I__7727\ : InMux
    port map (
            O => \N__37710\,
            I => \N__37700\
        );

    \I__7726\ : InMux
    port map (
            O => \N__37709\,
            I => \N__37697\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__37708\,
            I => \N__37694\
        );

    \I__7724\ : InMux
    port map (
            O => \N__37707\,
            I => \N__37689\
        );

    \I__7723\ : CascadeMux
    port map (
            O => \N__37706\,
            I => \N__37683\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__37703\,
            I => \N__37674\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__37700\,
            I => \N__37674\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__37697\,
            I => \N__37674\
        );

    \I__7719\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37660\
        );

    \I__7718\ : InMux
    port map (
            O => \N__37693\,
            I => \N__37655\
        );

    \I__7717\ : InMux
    port map (
            O => \N__37692\,
            I => \N__37655\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__37689\,
            I => \N__37652\
        );

    \I__7715\ : InMux
    port map (
            O => \N__37688\,
            I => \N__37643\
        );

    \I__7714\ : InMux
    port map (
            O => \N__37687\,
            I => \N__37643\
        );

    \I__7713\ : InMux
    port map (
            O => \N__37686\,
            I => \N__37643\
        );

    \I__7712\ : InMux
    port map (
            O => \N__37683\,
            I => \N__37643\
        );

    \I__7711\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37640\
        );

    \I__7710\ : InMux
    port map (
            O => \N__37681\,
            I => \N__37637\
        );

    \I__7709\ : Span4Mux_v
    port map (
            O => \N__37674\,
            I => \N__37634\
        );

    \I__7708\ : InMux
    port map (
            O => \N__37673\,
            I => \N__37631\
        );

    \I__7707\ : CascadeMux
    port map (
            O => \N__37672\,
            I => \N__37624\
        );

    \I__7706\ : CascadeMux
    port map (
            O => \N__37671\,
            I => \N__37621\
        );

    \I__7705\ : CascadeMux
    port map (
            O => \N__37670\,
            I => \N__37618\
        );

    \I__7704\ : CascadeMux
    port map (
            O => \N__37669\,
            I => \N__37615\
        );

    \I__7703\ : CascadeMux
    port map (
            O => \N__37668\,
            I => \N__37609\
        );

    \I__7702\ : CascadeMux
    port map (
            O => \N__37667\,
            I => \N__37606\
        );

    \I__7701\ : InMux
    port map (
            O => \N__37666\,
            I => \N__37603\
        );

    \I__7700\ : CascadeMux
    port map (
            O => \N__37665\,
            I => \N__37599\
        );

    \I__7699\ : InMux
    port map (
            O => \N__37664\,
            I => \N__37596\
        );

    \I__7698\ : InMux
    port map (
            O => \N__37663\,
            I => \N__37593\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__37660\,
            I => \N__37588\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__37655\,
            I => \N__37588\
        );

    \I__7695\ : Span4Mux_v
    port map (
            O => \N__37652\,
            I => \N__37583\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__37643\,
            I => \N__37583\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__37640\,
            I => \N__37578\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__37637\,
            I => \N__37578\
        );

    \I__7691\ : Span4Mux_h
    port map (
            O => \N__37634\,
            I => \N__37573\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__37631\,
            I => \N__37573\
        );

    \I__7689\ : InMux
    port map (
            O => \N__37630\,
            I => \N__37556\
        );

    \I__7688\ : InMux
    port map (
            O => \N__37629\,
            I => \N__37556\
        );

    \I__7687\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37556\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37627\,
            I => \N__37556\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37624\,
            I => \N__37556\
        );

    \I__7684\ : InMux
    port map (
            O => \N__37621\,
            I => \N__37556\
        );

    \I__7683\ : InMux
    port map (
            O => \N__37618\,
            I => \N__37556\
        );

    \I__7682\ : InMux
    port map (
            O => \N__37615\,
            I => \N__37556\
        );

    \I__7681\ : InMux
    port map (
            O => \N__37614\,
            I => \N__37545\
        );

    \I__7680\ : InMux
    port map (
            O => \N__37613\,
            I => \N__37545\
        );

    \I__7679\ : InMux
    port map (
            O => \N__37612\,
            I => \N__37545\
        );

    \I__7678\ : InMux
    port map (
            O => \N__37609\,
            I => \N__37545\
        );

    \I__7677\ : InMux
    port map (
            O => \N__37606\,
            I => \N__37545\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__37603\,
            I => \N__37542\
        );

    \I__7675\ : InMux
    port map (
            O => \N__37602\,
            I => \N__37537\
        );

    \I__7674\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37537\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__37596\,
            I => \N__37530\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__37593\,
            I => \N__37530\
        );

    \I__7671\ : Span4Mux_h
    port map (
            O => \N__37588\,
            I => \N__37530\
        );

    \I__7670\ : Span4Mux_h
    port map (
            O => \N__37583\,
            I => \N__37527\
        );

    \I__7669\ : Span12Mux_h
    port map (
            O => \N__37578\,
            I => \N__37524\
        );

    \I__7668\ : Span4Mux_h
    port map (
            O => \N__37573\,
            I => \N__37521\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__37556\,
            I => \N__37514\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__37545\,
            I => \N__37514\
        );

    \I__7665\ : Span12Mux_s7_v
    port map (
            O => \N__37542\,
            I => \N__37514\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__37537\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__37530\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__37527\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__7661\ : Odrv12
    port map (
            O => \N__37524\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__7660\ : Odrv4
    port map (
            O => \N__37521\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__7659\ : Odrv12
    port map (
            O => \N__37514\,
            I => \current_shift_inst.PI_CTRL.N_74\
        );

    \I__7658\ : InMux
    port map (
            O => \N__37501\,
            I => \N__37489\
        );

    \I__7657\ : InMux
    port map (
            O => \N__37500\,
            I => \N__37485\
        );

    \I__7656\ : InMux
    port map (
            O => \N__37499\,
            I => \N__37482\
        );

    \I__7655\ : InMux
    port map (
            O => \N__37498\,
            I => \N__37479\
        );

    \I__7654\ : InMux
    port map (
            O => \N__37497\,
            I => \N__37476\
        );

    \I__7653\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37464\
        );

    \I__7652\ : InMux
    port map (
            O => \N__37495\,
            I => \N__37464\
        );

    \I__7651\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37464\
        );

    \I__7650\ : InMux
    port map (
            O => \N__37493\,
            I => \N__37464\
        );

    \I__7649\ : InMux
    port map (
            O => \N__37492\,
            I => \N__37464\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__37489\,
            I => \N__37461\
        );

    \I__7647\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37457\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__37485\,
            I => \N__37435\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__37482\,
            I => \N__37432\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__37479\,
            I => \N__37427\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__37476\,
            I => \N__37427\
        );

    \I__7642\ : InMux
    port map (
            O => \N__37475\,
            I => \N__37424\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__37464\,
            I => \N__37419\
        );

    \I__7640\ : Span4Mux_h
    port map (
            O => \N__37461\,
            I => \N__37419\
        );

    \I__7639\ : InMux
    port map (
            O => \N__37460\,
            I => \N__37416\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__37457\,
            I => \N__37413\
        );

    \I__7637\ : InMux
    port map (
            O => \N__37456\,
            I => \N__37404\
        );

    \I__7636\ : InMux
    port map (
            O => \N__37455\,
            I => \N__37404\
        );

    \I__7635\ : InMux
    port map (
            O => \N__37454\,
            I => \N__37404\
        );

    \I__7634\ : InMux
    port map (
            O => \N__37453\,
            I => \N__37404\
        );

    \I__7633\ : InMux
    port map (
            O => \N__37452\,
            I => \N__37387\
        );

    \I__7632\ : InMux
    port map (
            O => \N__37451\,
            I => \N__37387\
        );

    \I__7631\ : InMux
    port map (
            O => \N__37450\,
            I => \N__37387\
        );

    \I__7630\ : InMux
    port map (
            O => \N__37449\,
            I => \N__37387\
        );

    \I__7629\ : InMux
    port map (
            O => \N__37448\,
            I => \N__37387\
        );

    \I__7628\ : InMux
    port map (
            O => \N__37447\,
            I => \N__37387\
        );

    \I__7627\ : InMux
    port map (
            O => \N__37446\,
            I => \N__37387\
        );

    \I__7626\ : InMux
    port map (
            O => \N__37445\,
            I => \N__37387\
        );

    \I__7625\ : InMux
    port map (
            O => \N__37444\,
            I => \N__37384\
        );

    \I__7624\ : InMux
    port map (
            O => \N__37443\,
            I => \N__37377\
        );

    \I__7623\ : InMux
    port map (
            O => \N__37442\,
            I => \N__37377\
        );

    \I__7622\ : InMux
    port map (
            O => \N__37441\,
            I => \N__37377\
        );

    \I__7621\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37372\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37372\
        );

    \I__7619\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37369\
        );

    \I__7618\ : Span4Mux_v
    port map (
            O => \N__37435\,
            I => \N__37366\
        );

    \I__7617\ : Span4Mux_v
    port map (
            O => \N__37432\,
            I => \N__37363\
        );

    \I__7616\ : Span12Mux_s9_v
    port map (
            O => \N__37427\,
            I => \N__37360\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__37424\,
            I => \N__37351\
        );

    \I__7614\ : Span4Mux_v
    port map (
            O => \N__37419\,
            I => \N__37351\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__37416\,
            I => \N__37351\
        );

    \I__7612\ : Span4Mux_v
    port map (
            O => \N__37413\,
            I => \N__37351\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__37404\,
            I => \N__37344\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__37387\,
            I => \N__37344\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__37384\,
            I => \N__37344\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__37377\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__37372\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__37369\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7605\ : Odrv4
    port map (
            O => \N__37366\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7604\ : Odrv4
    port map (
            O => \N__37363\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7603\ : Odrv12
    port map (
            O => \N__37360\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7602\ : Odrv4
    port map (
            O => \N__37351\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7601\ : Odrv4
    port map (
            O => \N__37344\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__7600\ : CascadeMux
    port map (
            O => \N__37327\,
            I => \N__37320\
        );

    \I__7599\ : CascadeMux
    port map (
            O => \N__37326\,
            I => \N__37317\
        );

    \I__7598\ : CascadeMux
    port map (
            O => \N__37325\,
            I => \N__37312\
        );

    \I__7597\ : CascadeMux
    port map (
            O => \N__37324\,
            I => \N__37309\
        );

    \I__7596\ : InMux
    port map (
            O => \N__37323\,
            I => \N__37304\
        );

    \I__7595\ : InMux
    port map (
            O => \N__37320\,
            I => \N__37300\
        );

    \I__7594\ : InMux
    port map (
            O => \N__37317\,
            I => \N__37297\
        );

    \I__7593\ : InMux
    port map (
            O => \N__37316\,
            I => \N__37294\
        );

    \I__7592\ : InMux
    port map (
            O => \N__37315\,
            I => \N__37291\
        );

    \I__7591\ : InMux
    port map (
            O => \N__37312\,
            I => \N__37277\
        );

    \I__7590\ : InMux
    port map (
            O => \N__37309\,
            I => \N__37277\
        );

    \I__7589\ : InMux
    port map (
            O => \N__37308\,
            I => \N__37274\
        );

    \I__7588\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37263\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__37304\,
            I => \N__37260\
        );

    \I__7586\ : InMux
    port map (
            O => \N__37303\,
            I => \N__37257\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__37300\,
            I => \N__37254\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__37297\,
            I => \N__37251\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__37294\,
            I => \N__37246\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__37291\,
            I => \N__37246\
        );

    \I__7581\ : InMux
    port map (
            O => \N__37290\,
            I => \N__37235\
        );

    \I__7580\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37235\
        );

    \I__7579\ : InMux
    port map (
            O => \N__37288\,
            I => \N__37235\
        );

    \I__7578\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37235\
        );

    \I__7577\ : InMux
    port map (
            O => \N__37286\,
            I => \N__37235\
        );

    \I__7576\ : InMux
    port map (
            O => \N__37285\,
            I => \N__37227\
        );

    \I__7575\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37224\
        );

    \I__7574\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37219\
        );

    \I__7573\ : InMux
    port map (
            O => \N__37282\,
            I => \N__37219\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__37277\,
            I => \N__37216\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__37274\,
            I => \N__37213\
        );

    \I__7570\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37196\
        );

    \I__7569\ : InMux
    port map (
            O => \N__37272\,
            I => \N__37196\
        );

    \I__7568\ : InMux
    port map (
            O => \N__37271\,
            I => \N__37196\
        );

    \I__7567\ : InMux
    port map (
            O => \N__37270\,
            I => \N__37196\
        );

    \I__7566\ : InMux
    port map (
            O => \N__37269\,
            I => \N__37196\
        );

    \I__7565\ : InMux
    port map (
            O => \N__37268\,
            I => \N__37196\
        );

    \I__7564\ : InMux
    port map (
            O => \N__37267\,
            I => \N__37196\
        );

    \I__7563\ : InMux
    port map (
            O => \N__37266\,
            I => \N__37196\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__37263\,
            I => \N__37191\
        );

    \I__7561\ : Span4Mux_h
    port map (
            O => \N__37260\,
            I => \N__37191\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__37257\,
            I => \N__37188\
        );

    \I__7559\ : Span4Mux_v
    port map (
            O => \N__37254\,
            I => \N__37183\
        );

    \I__7558\ : Span4Mux_v
    port map (
            O => \N__37251\,
            I => \N__37183\
        );

    \I__7557\ : Span4Mux_h
    port map (
            O => \N__37246\,
            I => \N__37178\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__37235\,
            I => \N__37178\
        );

    \I__7555\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37175\
        );

    \I__7554\ : InMux
    port map (
            O => \N__37233\,
            I => \N__37166\
        );

    \I__7553\ : InMux
    port map (
            O => \N__37232\,
            I => \N__37166\
        );

    \I__7552\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37166\
        );

    \I__7551\ : InMux
    port map (
            O => \N__37230\,
            I => \N__37166\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__37227\,
            I => \N__37161\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__37224\,
            I => \N__37161\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__37219\,
            I => \N__37158\
        );

    \I__7547\ : Span4Mux_v
    port map (
            O => \N__37216\,
            I => \N__37151\
        );

    \I__7546\ : Span4Mux_v
    port map (
            O => \N__37213\,
            I => \N__37151\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__37196\,
            I => \N__37151\
        );

    \I__7544\ : Span4Mux_h
    port map (
            O => \N__37191\,
            I => \N__37148\
        );

    \I__7543\ : Span4Mux_v
    port map (
            O => \N__37188\,
            I => \N__37143\
        );

    \I__7542\ : Span4Mux_h
    port map (
            O => \N__37183\,
            I => \N__37143\
        );

    \I__7541\ : Span4Mux_v
    port map (
            O => \N__37178\,
            I => \N__37140\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__37175\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__37166\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__7538\ : Odrv12
    port map (
            O => \N__37161\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__7537\ : Odrv12
    port map (
            O => \N__37158\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__7536\ : Odrv4
    port map (
            O => \N__37151\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__7535\ : Odrv4
    port map (
            O => \N__37148\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__37143\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__37140\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__7532\ : InMux
    port map (
            O => \N__37123\,
            I => \N__37120\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__37120\,
            I => \N__37117\
        );

    \I__7530\ : Odrv12
    port map (
            O => \N__37117\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__7529\ : CascadeMux
    port map (
            O => \N__37114\,
            I => \N__37111\
        );

    \I__7528\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37108\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__37108\,
            I => \N__37104\
        );

    \I__7526\ : InMux
    port map (
            O => \N__37107\,
            I => \N__37101\
        );

    \I__7525\ : Span4Mux_h
    port map (
            O => \N__37104\,
            I => \N__37095\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__37101\,
            I => \N__37095\
        );

    \I__7523\ : InMux
    port map (
            O => \N__37100\,
            I => \N__37092\
        );

    \I__7522\ : Span4Mux_v
    port map (
            O => \N__37095\,
            I => \N__37086\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__37092\,
            I => \N__37086\
        );

    \I__7520\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37083\
        );

    \I__7519\ : Span4Mux_h
    port map (
            O => \N__37086\,
            I => \N__37079\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__37083\,
            I => \N__37076\
        );

    \I__7517\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37073\
        );

    \I__7516\ : Span4Mux_h
    port map (
            O => \N__37079\,
            I => \N__37070\
        );

    \I__7515\ : Span4Mux_h
    port map (
            O => \N__37076\,
            I => \N__37067\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__37073\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__7513\ : Odrv4
    port map (
            O => \N__37070\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__7512\ : Odrv4
    port map (
            O => \N__37067\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__7511\ : InMux
    port map (
            O => \N__37060\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__7510\ : CascadeMux
    port map (
            O => \N__37057\,
            I => \N__37054\
        );

    \I__7509\ : InMux
    port map (
            O => \N__37054\,
            I => \N__37051\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__37051\,
            I => \N__37047\
        );

    \I__7507\ : InMux
    port map (
            O => \N__37050\,
            I => \N__37044\
        );

    \I__7506\ : Span4Mux_v
    port map (
            O => \N__37047\,
            I => \N__37037\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__37044\,
            I => \N__37037\
        );

    \I__7504\ : InMux
    port map (
            O => \N__37043\,
            I => \N__37034\
        );

    \I__7503\ : InMux
    port map (
            O => \N__37042\,
            I => \N__37031\
        );

    \I__7502\ : Sp12to4
    port map (
            O => \N__37037\,
            I => \N__37026\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__37034\,
            I => \N__37026\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__37031\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__7499\ : Odrv12
    port map (
            O => \N__37026\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__7498\ : InMux
    port map (
            O => \N__37021\,
            I => \N__37018\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__37018\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2\
        );

    \I__7496\ : InMux
    port map (
            O => \N__37015\,
            I => \N__37011\
        );

    \I__7495\ : InMux
    port map (
            O => \N__37014\,
            I => \N__37008\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__37011\,
            I => \N__37005\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__37008\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__7492\ : Odrv4
    port map (
            O => \N__37005\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__7491\ : InMux
    port map (
            O => \N__37000\,
            I => \N__36996\
        );

    \I__7490\ : InMux
    port map (
            O => \N__36999\,
            I => \N__36993\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__36996\,
            I => \N__36990\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__36993\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__36990\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__7486\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36982\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__36982\,
            I => \N__36979\
        );

    \I__7484\ : Span4Mux_h
    port map (
            O => \N__36979\,
            I => \N__36976\
        );

    \I__7483\ : Odrv4
    port map (
            O => \N__36976\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df20\
        );

    \I__7482\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36969\
        );

    \I__7481\ : InMux
    port map (
            O => \N__36972\,
            I => \N__36966\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__36969\,
            I => \N__36963\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__36966\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__36963\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36954\
        );

    \I__7476\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36951\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__36954\,
            I => \N__36948\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__36951\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__7473\ : Odrv4
    port map (
            O => \N__36948\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36943\,
            I => \N__36940\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__36940\,
            I => \N__36937\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__36937\,
            I => \N__36934\
        );

    \I__7469\ : Odrv4
    port map (
            O => \N__36934\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df22\
        );

    \I__7468\ : InMux
    port map (
            O => \N__36931\,
            I => \N__36927\
        );

    \I__7467\ : InMux
    port map (
            O => \N__36930\,
            I => \N__36924\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__36927\,
            I => \N__36921\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__36924\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__7464\ : Odrv4
    port map (
            O => \N__36921\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36916\,
            I => \N__36912\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36915\,
            I => \N__36909\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__36912\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__36909\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36904\,
            I => \N__36901\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36901\,
            I => \N__36898\
        );

    \I__7457\ : Span4Mux_v
    port map (
            O => \N__36898\,
            I => \N__36895\
        );

    \I__7456\ : Odrv4
    port map (
            O => \N__36895\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df24\
        );

    \I__7455\ : InMux
    port map (
            O => \N__36892\,
            I => \N__36888\
        );

    \I__7454\ : InMux
    port map (
            O => \N__36891\,
            I => \N__36885\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__36888\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__36885\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__7451\ : CascadeMux
    port map (
            O => \N__36880\,
            I => \N__36876\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36879\,
            I => \N__36873\
        );

    \I__7449\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36870\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__36873\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__36870\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__7446\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36862\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36859\
        );

    \I__7444\ : Span4Mux_v
    port map (
            O => \N__36859\,
            I => \N__36856\
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__36856\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df26\
        );

    \I__7442\ : InMux
    port map (
            O => \N__36853\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36850\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__7440\ : InMux
    port map (
            O => \N__36847\,
            I => \bfn_14_18_0_\
        );

    \I__7439\ : InMux
    port map (
            O => \N__36844\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__7438\ : InMux
    port map (
            O => \N__36841\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36838\,
            I => \N__36835\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36835\,
            I => \N__36831\
        );

    \I__7435\ : InMux
    port map (
            O => \N__36834\,
            I => \N__36828\
        );

    \I__7434\ : Span4Mux_v
    port map (
            O => \N__36831\,
            I => \N__36825\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__36828\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__7432\ : Odrv4
    port map (
            O => \N__36825\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36820\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__7430\ : InMux
    port map (
            O => \N__36817\,
            I => \N__36814\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__36814\,
            I => \N__36810\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36813\,
            I => \N__36807\
        );

    \I__7427\ : Span4Mux_v
    port map (
            O => \N__36810\,
            I => \N__36804\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__36807\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__36804\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36799\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__7423\ : InMux
    port map (
            O => \N__36796\,
            I => \N__36792\
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__36795\,
            I => \N__36789\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__36792\,
            I => \N__36785\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36789\,
            I => \N__36782\
        );

    \I__7419\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36779\
        );

    \I__7418\ : Span4Mux_v
    port map (
            O => \N__36785\,
            I => \N__36776\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__36782\,
            I => \N__36773\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__36779\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__7415\ : Odrv4
    port map (
            O => \N__36776\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__7414\ : Odrv12
    port map (
            O => \N__36773\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__7413\ : InMux
    port map (
            O => \N__36766\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__7412\ : CEMux
    port map (
            O => \N__36763\,
            I => \N__36758\
        );

    \I__7411\ : CEMux
    port map (
            O => \N__36762\,
            I => \N__36755\
        );

    \I__7410\ : CEMux
    port map (
            O => \N__36761\,
            I => \N__36751\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__36758\,
            I => \N__36740\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__36755\,
            I => \N__36736\
        );

    \I__7407\ : CEMux
    port map (
            O => \N__36754\,
            I => \N__36733\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__36751\,
            I => \N__36730\
        );

    \I__7405\ : CEMux
    port map (
            O => \N__36750\,
            I => \N__36716\
        );

    \I__7404\ : InMux
    port map (
            O => \N__36749\,
            I => \N__36709\
        );

    \I__7403\ : InMux
    port map (
            O => \N__36748\,
            I => \N__36709\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36747\,
            I => \N__36709\
        );

    \I__7401\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36700\
        );

    \I__7400\ : InMux
    port map (
            O => \N__36745\,
            I => \N__36700\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36744\,
            I => \N__36700\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36700\
        );

    \I__7397\ : Span4Mux_v
    port map (
            O => \N__36740\,
            I => \N__36685\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36739\,
            I => \N__36682\
        );

    \I__7395\ : Span4Mux_v
    port map (
            O => \N__36736\,
            I => \N__36677\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__36733\,
            I => \N__36677\
        );

    \I__7393\ : Span4Mux_h
    port map (
            O => \N__36730\,
            I => \N__36674\
        );

    \I__7392\ : InMux
    port map (
            O => \N__36729\,
            I => \N__36665\
        );

    \I__7391\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36665\
        );

    \I__7390\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36665\
        );

    \I__7389\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36665\
        );

    \I__7388\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36656\
        );

    \I__7387\ : InMux
    port map (
            O => \N__36724\,
            I => \N__36656\
        );

    \I__7386\ : InMux
    port map (
            O => \N__36723\,
            I => \N__36656\
        );

    \I__7385\ : InMux
    port map (
            O => \N__36722\,
            I => \N__36656\
        );

    \I__7384\ : InMux
    port map (
            O => \N__36721\,
            I => \N__36649\
        );

    \I__7383\ : InMux
    port map (
            O => \N__36720\,
            I => \N__36649\
        );

    \I__7382\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36649\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__36716\,
            I => \N__36646\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__36709\,
            I => \N__36641\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__36700\,
            I => \N__36641\
        );

    \I__7378\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36632\
        );

    \I__7377\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36632\
        );

    \I__7376\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36632\
        );

    \I__7375\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36632\
        );

    \I__7374\ : InMux
    port map (
            O => \N__36695\,
            I => \N__36623\
        );

    \I__7373\ : InMux
    port map (
            O => \N__36694\,
            I => \N__36623\
        );

    \I__7372\ : InMux
    port map (
            O => \N__36693\,
            I => \N__36623\
        );

    \I__7371\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36623\
        );

    \I__7370\ : InMux
    port map (
            O => \N__36691\,
            I => \N__36614\
        );

    \I__7369\ : InMux
    port map (
            O => \N__36690\,
            I => \N__36614\
        );

    \I__7368\ : InMux
    port map (
            O => \N__36689\,
            I => \N__36614\
        );

    \I__7367\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36614\
        );

    \I__7366\ : Span4Mux_h
    port map (
            O => \N__36685\,
            I => \N__36609\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__36682\,
            I => \N__36609\
        );

    \I__7364\ : Span4Mux_v
    port map (
            O => \N__36677\,
            I => \N__36606\
        );

    \I__7363\ : Span4Mux_v
    port map (
            O => \N__36674\,
            I => \N__36601\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__36665\,
            I => \N__36601\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__36656\,
            I => \N__36598\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__36649\,
            I => \N__36585\
        );

    \I__7359\ : Span4Mux_v
    port map (
            O => \N__36646\,
            I => \N__36585\
        );

    \I__7358\ : Span4Mux_h
    port map (
            O => \N__36641\,
            I => \N__36585\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__36632\,
            I => \N__36585\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__36623\,
            I => \N__36585\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__36614\,
            I => \N__36585\
        );

    \I__7354\ : Span4Mux_v
    port map (
            O => \N__36609\,
            I => \N__36582\
        );

    \I__7353\ : Span4Mux_h
    port map (
            O => \N__36606\,
            I => \N__36579\
        );

    \I__7352\ : Span4Mux_h
    port map (
            O => \N__36601\,
            I => \N__36576\
        );

    \I__7351\ : Span4Mux_v
    port map (
            O => \N__36598\,
            I => \N__36571\
        );

    \I__7350\ : Span4Mux_v
    port map (
            O => \N__36585\,
            I => \N__36571\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__36582\,
            I => \N__36568\
        );

    \I__7348\ : Span4Mux_v
    port map (
            O => \N__36579\,
            I => \N__36565\
        );

    \I__7347\ : Odrv4
    port map (
            O => \N__36576\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__7346\ : Odrv4
    port map (
            O => \N__36571\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__36568\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__36565\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__7343\ : InMux
    port map (
            O => \N__36556\,
            I => \N__36552\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36555\,
            I => \N__36549\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__36552\,
            I => \N__36546\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__36549\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__36546\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7338\ : InMux
    port map (
            O => \N__36541\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__7337\ : InMux
    port map (
            O => \N__36538\,
            I => \N__36535\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__36535\,
            I => \N__36531\
        );

    \I__7335\ : InMux
    port map (
            O => \N__36534\,
            I => \N__36528\
        );

    \I__7334\ : Span4Mux_v
    port map (
            O => \N__36531\,
            I => \N__36525\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__36528\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7332\ : Odrv4
    port map (
            O => \N__36525\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7331\ : InMux
    port map (
            O => \N__36520\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__7330\ : CascadeMux
    port map (
            O => \N__36517\,
            I => \N__36513\
        );

    \I__7329\ : CascadeMux
    port map (
            O => \N__36516\,
            I => \N__36510\
        );

    \I__7328\ : InMux
    port map (
            O => \N__36513\,
            I => \N__36507\
        );

    \I__7327\ : InMux
    port map (
            O => \N__36510\,
            I => \N__36504\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__36507\,
            I => \N__36501\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__36504\,
            I => \N__36497\
        );

    \I__7324\ : Span4Mux_h
    port map (
            O => \N__36501\,
            I => \N__36494\
        );

    \I__7323\ : InMux
    port map (
            O => \N__36500\,
            I => \N__36491\
        );

    \I__7322\ : Span4Mux_v
    port map (
            O => \N__36497\,
            I => \N__36486\
        );

    \I__7321\ : Span4Mux_v
    port map (
            O => \N__36494\,
            I => \N__36486\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__36491\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__7319\ : Odrv4
    port map (
            O => \N__36486\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__7318\ : InMux
    port map (
            O => \N__36481\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__7317\ : InMux
    port map (
            O => \N__36478\,
            I => \N__36474\
        );

    \I__7316\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36470\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__36474\,
            I => \N__36467\
        );

    \I__7314\ : InMux
    port map (
            O => \N__36473\,
            I => \N__36464\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__36470\,
            I => \N__36461\
        );

    \I__7312\ : Span4Mux_h
    port map (
            O => \N__36467\,
            I => \N__36458\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__36464\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7310\ : Odrv12
    port map (
            O => \N__36461\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7309\ : Odrv4
    port map (
            O => \N__36458\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7308\ : InMux
    port map (
            O => \N__36451\,
            I => \bfn_14_17_0_\
        );

    \I__7307\ : CascadeMux
    port map (
            O => \N__36448\,
            I => \N__36444\
        );

    \I__7306\ : InMux
    port map (
            O => \N__36447\,
            I => \N__36439\
        );

    \I__7305\ : InMux
    port map (
            O => \N__36444\,
            I => \N__36439\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__36439\,
            I => \N__36435\
        );

    \I__7303\ : InMux
    port map (
            O => \N__36438\,
            I => \N__36432\
        );

    \I__7302\ : Span4Mux_v
    port map (
            O => \N__36435\,
            I => \N__36429\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__36432\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__36429\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__7299\ : InMux
    port map (
            O => \N__36424\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__7298\ : InMux
    port map (
            O => \N__36421\,
            I => \N__36414\
        );

    \I__7297\ : InMux
    port map (
            O => \N__36420\,
            I => \N__36414\
        );

    \I__7296\ : InMux
    port map (
            O => \N__36419\,
            I => \N__36411\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__36414\,
            I => \N__36408\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__36411\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7293\ : Odrv12
    port map (
            O => \N__36408\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__7292\ : InMux
    port map (
            O => \N__36403\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__7291\ : InMux
    port map (
            O => \N__36400\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__7290\ : InMux
    port map (
            O => \N__36397\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__7289\ : InMux
    port map (
            O => \N__36394\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__7288\ : InMux
    port map (
            O => \N__36391\,
            I => \N__36388\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__36388\,
            I => \N__36384\
        );

    \I__7286\ : InMux
    port map (
            O => \N__36387\,
            I => \N__36381\
        );

    \I__7285\ : Span4Mux_h
    port map (
            O => \N__36384\,
            I => \N__36378\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__36381\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7283\ : Odrv4
    port map (
            O => \N__36378\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7282\ : InMux
    port map (
            O => \N__36373\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__7281\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36366\
        );

    \I__7280\ : InMux
    port map (
            O => \N__36369\,
            I => \N__36363\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__36366\,
            I => \N__36360\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__36363\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7277\ : Odrv4
    port map (
            O => \N__36360\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7276\ : InMux
    port map (
            O => \N__36355\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__7275\ : InMux
    port map (
            O => \N__36352\,
            I => \N__36348\
        );

    \I__7274\ : InMux
    port map (
            O => \N__36351\,
            I => \N__36345\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__36348\,
            I => \N__36342\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__36345\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7271\ : Odrv4
    port map (
            O => \N__36342\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36337\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__7269\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36330\
        );

    \I__7268\ : InMux
    port map (
            O => \N__36333\,
            I => \N__36327\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__36330\,
            I => \N__36324\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__36327\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7265\ : Odrv4
    port map (
            O => \N__36324\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7264\ : InMux
    port map (
            O => \N__36319\,
            I => \bfn_14_16_0_\
        );

    \I__7263\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36312\
        );

    \I__7262\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36309\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__36312\,
            I => \N__36306\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__36309\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7259\ : Odrv4
    port map (
            O => \N__36306\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7258\ : InMux
    port map (
            O => \N__36301\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__7257\ : InMux
    port map (
            O => \N__36298\,
            I => \N__36295\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__36295\,
            I => \N__36292\
        );

    \I__7255\ : Span4Mux_v
    port map (
            O => \N__36292\,
            I => \N__36288\
        );

    \I__7254\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36285\
        );

    \I__7253\ : Sp12to4
    port map (
            O => \N__36288\,
            I => \N__36282\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__36285\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7251\ : Odrv12
    port map (
            O => \N__36282\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7250\ : InMux
    port map (
            O => \N__36277\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__7249\ : InMux
    port map (
            O => \N__36274\,
            I => \N__36270\
        );

    \I__7248\ : InMux
    port map (
            O => \N__36273\,
            I => \N__36267\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__36270\,
            I => \N__36264\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__36267\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7245\ : Odrv4
    port map (
            O => \N__36264\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7244\ : InMux
    port map (
            O => \N__36259\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__7243\ : InMux
    port map (
            O => \N__36256\,
            I => \N__36252\
        );

    \I__7242\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36249\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__36252\,
            I => \N__36246\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__36249\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7239\ : Odrv4
    port map (
            O => \N__36246\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7238\ : InMux
    port map (
            O => \N__36241\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__7237\ : InMux
    port map (
            O => \N__36238\,
            I => \N__36235\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__36235\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__7235\ : CascadeMux
    port map (
            O => \N__36232\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__7234\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36225\
        );

    \I__7233\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36219\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__36225\,
            I => \N__36216\
        );

    \I__7231\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36209\
        );

    \I__7230\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36209\
        );

    \I__7229\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36209\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__36219\,
            I => \N__36206\
        );

    \I__7227\ : Span4Mux_v
    port map (
            O => \N__36216\,
            I => \N__36201\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__36209\,
            I => \N__36201\
        );

    \I__7225\ : Span4Mux_v
    port map (
            O => \N__36206\,
            I => \N__36198\
        );

    \I__7224\ : Span4Mux_h
    port map (
            O => \N__36201\,
            I => \N__36195\
        );

    \I__7223\ : Odrv4
    port map (
            O => \N__36198\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__7222\ : Odrv4
    port map (
            O => \N__36195\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__7221\ : InMux
    port map (
            O => \N__36190\,
            I => \N__36184\
        );

    \I__7220\ : InMux
    port map (
            O => \N__36189\,
            I => \N__36184\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__36184\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__7218\ : InMux
    port map (
            O => \N__36181\,
            I => \N__36177\
        );

    \I__7217\ : InMux
    port map (
            O => \N__36180\,
            I => \N__36174\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__36177\,
            I => \N__36171\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__36174\,
            I => \N__36167\
        );

    \I__7214\ : Span4Mux_v
    port map (
            O => \N__36171\,
            I => \N__36164\
        );

    \I__7213\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36160\
        );

    \I__7212\ : Span4Mux_h
    port map (
            O => \N__36167\,
            I => \N__36157\
        );

    \I__7211\ : Span4Mux_h
    port map (
            O => \N__36164\,
            I => \N__36154\
        );

    \I__7210\ : InMux
    port map (
            O => \N__36163\,
            I => \N__36151\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__36160\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7208\ : Odrv4
    port map (
            O => \N__36157\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__36154\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__36151\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7205\ : CascadeMux
    port map (
            O => \N__36142\,
            I => \N__36137\
        );

    \I__7204\ : InMux
    port map (
            O => \N__36141\,
            I => \N__36132\
        );

    \I__7203\ : InMux
    port map (
            O => \N__36140\,
            I => \N__36132\
        );

    \I__7202\ : InMux
    port map (
            O => \N__36137\,
            I => \N__36129\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__36132\,
            I => \N__36126\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__36129\,
            I => \N__36122\
        );

    \I__7199\ : Span4Mux_h
    port map (
            O => \N__36126\,
            I => \N__36119\
        );

    \I__7198\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36116\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__36122\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__7196\ : Odrv4
    port map (
            O => \N__36119\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__36116\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__7194\ : CascadeMux
    port map (
            O => \N__36109\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\
        );

    \I__7193\ : InMux
    port map (
            O => \N__36106\,
            I => \N__36103\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__36103\,
            I => \N__36100\
        );

    \I__7191\ : Span4Mux_h
    port map (
            O => \N__36100\,
            I => \N__36096\
        );

    \I__7190\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36093\
        );

    \I__7189\ : Odrv4
    port map (
            O => \N__36096\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__36093\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__7187\ : InMux
    port map (
            O => \N__36088\,
            I => \N__36085\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__36085\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__7185\ : CascadeMux
    port map (
            O => \N__36082\,
            I => \N__36079\
        );

    \I__7184\ : InMux
    port map (
            O => \N__36079\,
            I => \N__36075\
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__36078\,
            I => \N__36071\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__36075\,
            I => \N__36068\
        );

    \I__7181\ : InMux
    port map (
            O => \N__36074\,
            I => \N__36065\
        );

    \I__7180\ : InMux
    port map (
            O => \N__36071\,
            I => \N__36062\
        );

    \I__7179\ : Span4Mux_h
    port map (
            O => \N__36068\,
            I => \N__36059\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__36065\,
            I => \N__36056\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__36062\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7176\ : Odrv4
    port map (
            O => \N__36059\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7175\ : Odrv4
    port map (
            O => \N__36056\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7174\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36045\
        );

    \I__7173\ : InMux
    port map (
            O => \N__36048\,
            I => \N__36042\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__36045\,
            I => \N__36039\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__36042\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7170\ : Odrv4
    port map (
            O => \N__36039\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7169\ : InMux
    port map (
            O => \N__36034\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__7168\ : CascadeMux
    port map (
            O => \N__36031\,
            I => \N__36028\
        );

    \I__7167\ : InMux
    port map (
            O => \N__36028\,
            I => \N__36025\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__36025\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28\
        );

    \I__7165\ : InMux
    port map (
            O => \N__36022\,
            I => \N__36018\
        );

    \I__7164\ : InMux
    port map (
            O => \N__36021\,
            I => \N__36015\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__36018\,
            I => \N__36012\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__36015\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__36012\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7160\ : InMux
    port map (
            O => \N__36007\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__7159\ : InMux
    port map (
            O => \N__36004\,
            I => \N__36000\
        );

    \I__7158\ : InMux
    port map (
            O => \N__36003\,
            I => \N__35997\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__36000\,
            I => \N__35994\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__35997\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7155\ : Odrv4
    port map (
            O => \N__35994\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35989\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__7153\ : InMux
    port map (
            O => \N__35986\,
            I => \N__35982\
        );

    \I__7152\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35979\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__35982\,
            I => \N__35976\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35979\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7149\ : Odrv4
    port map (
            O => \N__35976\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35971\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__7147\ : CascadeMux
    port map (
            O => \N__35968\,
            I => \N__35965\
        );

    \I__7146\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35962\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__35962\,
            I => \N__35959\
        );

    \I__7144\ : Span4Mux_v
    port map (
            O => \N__35959\,
            I => \N__35956\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__35956\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__7142\ : CascadeMux
    port map (
            O => \N__35953\,
            I => \N__35950\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35944\
        );

    \I__7140\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35944\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__35944\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__7138\ : InMux
    port map (
            O => \N__35941\,
            I => \N__35938\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__35938\,
            I => \N__35935\
        );

    \I__7136\ : Odrv4
    port map (
            O => \N__35935\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__7135\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35926\
        );

    \I__7134\ : InMux
    port map (
            O => \N__35931\,
            I => \N__35926\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__35926\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35923\,
            I => \N__35919\
        );

    \I__7131\ : InMux
    port map (
            O => \N__35922\,
            I => \N__35916\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35919\,
            I => \N__35913\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__35916\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__7128\ : Odrv12
    port map (
            O => \N__35913\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35908\,
            I => \N__35905\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__35905\,
            I => \N__35901\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35904\,
            I => \N__35898\
        );

    \I__7124\ : Span4Mux_v
    port map (
            O => \N__35901\,
            I => \N__35895\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__35898\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__7122\ : Odrv4
    port map (
            O => \N__35895\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__7121\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35887\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__35887\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__7119\ : InMux
    port map (
            O => \N__35884\,
            I => \N__35880\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35883\,
            I => \N__35877\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35880\,
            I => \N__35874\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__35877\,
            I => \N__35869\
        );

    \I__7115\ : Span12Mux_h
    port map (
            O => \N__35874\,
            I => \N__35866\
        );

    \I__7114\ : InMux
    port map (
            O => \N__35873\,
            I => \N__35863\
        );

    \I__7113\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35860\
        );

    \I__7112\ : Span4Mux_h
    port map (
            O => \N__35869\,
            I => \N__35857\
        );

    \I__7111\ : Span12Mux_v
    port map (
            O => \N__35866\,
            I => \N__35854\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35863\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__35860\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__7108\ : Odrv4
    port map (
            O => \N__35857\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__7107\ : Odrv12
    port map (
            O => \N__35854\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__7106\ : InMux
    port map (
            O => \N__35845\,
            I => \N__35838\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35838\
        );

    \I__7104\ : InMux
    port map (
            O => \N__35843\,
            I => \N__35835\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__35838\,
            I => \N__35832\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__35835\,
            I => \N__35829\
        );

    \I__7101\ : Span4Mux_v
    port map (
            O => \N__35832\,
            I => \N__35824\
        );

    \I__7100\ : Span4Mux_h
    port map (
            O => \N__35829\,
            I => \N__35824\
        );

    \I__7099\ : Span4Mux_h
    port map (
            O => \N__35824\,
            I => \N__35821\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__35821\,
            I => \il_min_comp2_D2\
        );

    \I__7097\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35814\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35811\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35808\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__35811\,
            I => \N__35803\
        );

    \I__7093\ : Span4Mux_v
    port map (
            O => \N__35808\,
            I => \N__35803\
        );

    \I__7092\ : Span4Mux_v
    port map (
            O => \N__35803\,
            I => \N__35800\
        );

    \I__7091\ : Odrv4
    port map (
            O => \N__35800\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__7090\ : CascadeMux
    port map (
            O => \N__35797\,
            I => \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_\
        );

    \I__7089\ : InMux
    port map (
            O => \N__35794\,
            I => \N__35790\
        );

    \I__7088\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35787\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__35790\,
            I => \N__35784\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__35787\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__7085\ : Odrv4
    port map (
            O => \N__35784\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__7084\ : CascadeMux
    port map (
            O => \N__35779\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35776\,
            I => \N__35773\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__35773\,
            I => \N__35769\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35772\,
            I => \N__35766\
        );

    \I__7080\ : Odrv4
    port map (
            O => \N__35769\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__35766\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2\
        );

    \I__7078\ : CascadeMux
    port map (
            O => \N__35761\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__35758\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_\
        );

    \I__7076\ : CascadeMux
    port map (
            O => \N__35755\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_\
        );

    \I__7075\ : InMux
    port map (
            O => \N__35752\,
            I => \N__35749\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__35749\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35746\,
            I => \N__35743\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__35743\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__7071\ : InMux
    port map (
            O => \N__35740\,
            I => \N__35737\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__35737\,
            I => \N__35734\
        );

    \I__7069\ : Span4Mux_h
    port map (
            O => \N__35734\,
            I => \N__35730\
        );

    \I__7068\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35727\
        );

    \I__7067\ : Odrv4
    port map (
            O => \N__35730\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__35727\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\
        );

    \I__7065\ : CascadeMux
    port map (
            O => \N__35722\,
            I => \elapsed_time_ns_1_RNIP7HF91_0_10_cascade_\
        );

    \I__7064\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35716\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__35716\,
            I => \N__35711\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35715\,
            I => \N__35708\
        );

    \I__7061\ : InMux
    port map (
            O => \N__35714\,
            I => \N__35704\
        );

    \I__7060\ : Span4Mux_v
    port map (
            O => \N__35711\,
            I => \N__35701\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__35708\,
            I => \N__35698\
        );

    \I__7058\ : InMux
    port map (
            O => \N__35707\,
            I => \N__35695\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__35704\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__7056\ : Odrv4
    port map (
            O => \N__35701\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__35698\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__35695\,
            I => \elapsed_time_ns_1_RNIFJ2591_0_7\
        );

    \I__7053\ : CascadeMux
    port map (
            O => \N__35686\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_\
        );

    \I__7052\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35680\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__35680\,
            I => \N__35677\
        );

    \I__7050\ : Span4Mux_v
    port map (
            O => \N__35677\,
            I => \N__35671\
        );

    \I__7049\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35668\
        );

    \I__7048\ : InMux
    port map (
            O => \N__35675\,
            I => \N__35663\
        );

    \I__7047\ : InMux
    port map (
            O => \N__35674\,
            I => \N__35663\
        );

    \I__7046\ : Odrv4
    port map (
            O => \N__35671\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__35668\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__35663\,
            I => \elapsed_time_ns_1_RNIGK2591_0_8\
        );

    \I__7043\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35652\
        );

    \I__7042\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35647\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__35652\,
            I => \N__35644\
        );

    \I__7040\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35641\
        );

    \I__7039\ : InMux
    port map (
            O => \N__35650\,
            I => \N__35638\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__35647\,
            I => \N__35635\
        );

    \I__7037\ : Span4Mux_h
    port map (
            O => \N__35644\,
            I => \N__35629\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__35641\,
            I => \N__35629\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__35638\,
            I => \N__35626\
        );

    \I__7034\ : Span4Mux_v
    port map (
            O => \N__35635\,
            I => \N__35623\
        );

    \I__7033\ : InMux
    port map (
            O => \N__35634\,
            I => \N__35620\
        );

    \I__7032\ : Span4Mux_h
    port map (
            O => \N__35629\,
            I => \N__35617\
        );

    \I__7031\ : Odrv12
    port map (
            O => \N__35626\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7030\ : Odrv4
    port map (
            O => \N__35623\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__35620\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7028\ : Odrv4
    port map (
            O => \N__35617\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7027\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35605\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__35605\,
            I => \N__35602\
        );

    \I__7025\ : Odrv12
    port map (
            O => \N__35602\,
            I => \current_shift_inst.PI_CTRL.integrator_i_19\
        );

    \I__7024\ : InMux
    port map (
            O => \N__35599\,
            I => \N__35596\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__35596\,
            I => \N__35593\
        );

    \I__7022\ : Span4Mux_h
    port map (
            O => \N__35593\,
            I => \N__35590\
        );

    \I__7021\ : Odrv4
    port map (
            O => \N__35590\,
            I => \current_shift_inst.PI_CTRL.integrator_i_9\
        );

    \I__7020\ : CascadeMux
    port map (
            O => \N__35587\,
            I => \N__35584\
        );

    \I__7019\ : InMux
    port map (
            O => \N__35584\,
            I => \N__35580\
        );

    \I__7018\ : InMux
    port map (
            O => \N__35583\,
            I => \N__35576\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__35580\,
            I => \N__35573\
        );

    \I__7016\ : InMux
    port map (
            O => \N__35579\,
            I => \N__35570\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__35576\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__35573\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__35570\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\
        );

    \I__7012\ : CascadeMux
    port map (
            O => \N__35563\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9_cascade_\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__35560\,
            I => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\
        );

    \I__7010\ : CascadeMux
    port map (
            O => \N__35557\,
            I => \N__35554\
        );

    \I__7009\ : InMux
    port map (
            O => \N__35554\,
            I => \N__35551\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__35551\,
            I => \N__35548\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__35548\,
            I => \N__35545\
        );

    \I__7006\ : Odrv4
    port map (
            O => \N__35545\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__7005\ : InMux
    port map (
            O => \N__35542\,
            I => \N__35539\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__35539\,
            I => \N__35536\
        );

    \I__7003\ : Span4Mux_v
    port map (
            O => \N__35536\,
            I => \N__35533\
        );

    \I__7002\ : Odrv4
    port map (
            O => \N__35533\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__35530\,
            I => \N__35527\
        );

    \I__7000\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35524\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__35524\,
            I => \N__35521\
        );

    \I__6998\ : Span4Mux_v
    port map (
            O => \N__35521\,
            I => \N__35518\
        );

    \I__6997\ : Odrv4
    port map (
            O => \N__35518\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__6996\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35511\
        );

    \I__6995\ : InMux
    port map (
            O => \N__35514\,
            I => \N__35507\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__35511\,
            I => \N__35504\
        );

    \I__6993\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35501\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__35507\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__6991\ : Odrv4
    port map (
            O => \N__35504\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__35501\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\
        );

    \I__6989\ : CascadeMux
    port map (
            O => \N__35494\,
            I => \N__35491\
        );

    \I__6988\ : InMux
    port map (
            O => \N__35491\,
            I => \N__35487\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35490\,
            I => \N__35483\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__35487\,
            I => \N__35480\
        );

    \I__6985\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35477\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__35483\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__6983\ : Odrv4
    port map (
            O => \N__35480\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__35477\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\
        );

    \I__6981\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35466\
        );

    \I__6980\ : InMux
    port map (
            O => \N__35469\,
            I => \N__35463\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__35466\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__35463\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\
        );

    \I__6977\ : InMux
    port map (
            O => \N__35458\,
            I => \N__35453\
        );

    \I__6976\ : InMux
    port map (
            O => \N__35457\,
            I => \N__35450\
        );

    \I__6975\ : InMux
    port map (
            O => \N__35456\,
            I => \N__35447\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__35453\,
            I => \N__35443\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__35450\,
            I => \N__35439\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__35447\,
            I => \N__35436\
        );

    \I__6971\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35433\
        );

    \I__6970\ : Span4Mux_v
    port map (
            O => \N__35443\,
            I => \N__35430\
        );

    \I__6969\ : InMux
    port map (
            O => \N__35442\,
            I => \N__35427\
        );

    \I__6968\ : Span4Mux_h
    port map (
            O => \N__35439\,
            I => \N__35422\
        );

    \I__6967\ : Span4Mux_h
    port map (
            O => \N__35436\,
            I => \N__35422\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__35433\,
            I => \N__35419\
        );

    \I__6965\ : Sp12to4
    port map (
            O => \N__35430\,
            I => \N__35414\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__35427\,
            I => \N__35414\
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__35422\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__6962\ : Odrv12
    port map (
            O => \N__35419\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__6961\ : Odrv12
    port map (
            O => \N__35414\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__35407\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28_cascade_\
        );

    \I__6959\ : InMux
    port map (
            O => \N__35404\,
            I => \N__35401\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__35401\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\
        );

    \I__6957\ : CascadeMux
    port map (
            O => \N__35398\,
            I => \N__35395\
        );

    \I__6956\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35392\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__35392\,
            I => \N__35389\
        );

    \I__6954\ : Span4Mux_h
    port map (
            O => \N__35389\,
            I => \N__35386\
        );

    \I__6953\ : Odrv4
    port map (
            O => \N__35386\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0\
        );

    \I__6952\ : InMux
    port map (
            O => \N__35383\,
            I => \N__35379\
        );

    \I__6951\ : InMux
    port map (
            O => \N__35382\,
            I => \N__35376\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__35379\,
            I => \N__35373\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__35376\,
            I => \N__35370\
        );

    \I__6948\ : Span4Mux_h
    port map (
            O => \N__35373\,
            I => \N__35367\
        );

    \I__6947\ : Span4Mux_v
    port map (
            O => \N__35370\,
            I => \N__35362\
        );

    \I__6946\ : Span4Mux_v
    port map (
            O => \N__35367\,
            I => \N__35359\
        );

    \I__6945\ : InMux
    port map (
            O => \N__35366\,
            I => \N__35356\
        );

    \I__6944\ : InMux
    port map (
            O => \N__35365\,
            I => \N__35353\
        );

    \I__6943\ : Span4Mux_h
    port map (
            O => \N__35362\,
            I => \N__35348\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__35359\,
            I => \N__35348\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__35356\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__35353\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6939\ : Odrv4
    port map (
            O => \N__35348\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6938\ : InMux
    port map (
            O => \N__35341\,
            I => \N__35336\
        );

    \I__6937\ : InMux
    port map (
            O => \N__35340\,
            I => \N__35333\
        );

    \I__6936\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35330\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__35336\,
            I => \N__35327\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__35333\,
            I => \N__35324\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__35330\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__6932\ : Odrv4
    port map (
            O => \N__35327\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__6931\ : Odrv4
    port map (
            O => \N__35324\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\
        );

    \I__6930\ : InMux
    port map (
            O => \N__35317\,
            I => \N__35314\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__35314\,
            I => \N__35311\
        );

    \I__6928\ : Odrv12
    port map (
            O => \N__35311\,
            I => \current_shift_inst.PI_CTRL.integrator_i_16\
        );

    \I__6927\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35303\
        );

    \I__6926\ : CascadeMux
    port map (
            O => \N__35307\,
            I => \N__35300\
        );

    \I__6925\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35297\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__35303\,
            I => \N__35294\
        );

    \I__6923\ : InMux
    port map (
            O => \N__35300\,
            I => \N__35291\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__35297\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__35294\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__35291\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\
        );

    \I__6919\ : CascadeMux
    port map (
            O => \N__35284\,
            I => \N__35280\
        );

    \I__6918\ : InMux
    port map (
            O => \N__35283\,
            I => \N__35277\
        );

    \I__6917\ : InMux
    port map (
            O => \N__35280\,
            I => \N__35274\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__35277\,
            I => \N__35270\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__35274\,
            I => \N__35267\
        );

    \I__6914\ : InMux
    port map (
            O => \N__35273\,
            I => \N__35262\
        );

    \I__6913\ : Span4Mux_v
    port map (
            O => \N__35270\,
            I => \N__35259\
        );

    \I__6912\ : Span4Mux_v
    port map (
            O => \N__35267\,
            I => \N__35256\
        );

    \I__6911\ : InMux
    port map (
            O => \N__35266\,
            I => \N__35251\
        );

    \I__6910\ : InMux
    port map (
            O => \N__35265\,
            I => \N__35251\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__35262\,
            I => \N__35248\
        );

    \I__6908\ : Odrv4
    port map (
            O => \N__35259\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__35256\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__35251\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__6905\ : Odrv4
    port map (
            O => \N__35248\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__6904\ : CascadeMux
    port map (
            O => \N__35239\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_\
        );

    \I__6903\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35233\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__35233\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__35230\,
            I => \N__35227\
        );

    \I__6900\ : InMux
    port map (
            O => \N__35227\,
            I => \N__35224\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__35224\,
            I => \N__35221\
        );

    \I__6898\ : Span12Mux_h
    port map (
            O => \N__35221\,
            I => \N__35218\
        );

    \I__6897\ : Odrv12
    port map (
            O => \N__35218\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0\
        );

    \I__6896\ : InMux
    port map (
            O => \N__35215\,
            I => \N__35212\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__35212\,
            I => \N__35208\
        );

    \I__6894\ : InMux
    port map (
            O => \N__35211\,
            I => \N__35204\
        );

    \I__6893\ : Span4Mux_h
    port map (
            O => \N__35208\,
            I => \N__35201\
        );

    \I__6892\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35198\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__35204\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__35201\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__35198\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\
        );

    \I__6888\ : CascadeMux
    port map (
            O => \N__35191\,
            I => \N__35187\
        );

    \I__6887\ : InMux
    port map (
            O => \N__35190\,
            I => \N__35184\
        );

    \I__6886\ : InMux
    port map (
            O => \N__35187\,
            I => \N__35180\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__35184\,
            I => \N__35177\
        );

    \I__6884\ : InMux
    port map (
            O => \N__35183\,
            I => \N__35174\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__35180\,
            I => \N__35171\
        );

    \I__6882\ : Span4Mux_h
    port map (
            O => \N__35177\,
            I => \N__35168\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__35174\,
            I => \N__35165\
        );

    \I__6880\ : Span4Mux_h
    port map (
            O => \N__35171\,
            I => \N__35162\
        );

    \I__6879\ : Span4Mux_v
    port map (
            O => \N__35168\,
            I => \N__35159\
        );

    \I__6878\ : Odrv4
    port map (
            O => \N__35165\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__35162\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6876\ : Odrv4
    port map (
            O => \N__35159\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__6875\ : InMux
    port map (
            O => \N__35152\,
            I => \N__35149\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__35149\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_12\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__35146\,
            I => \N__35143\
        );

    \I__6872\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35140\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__35140\,
            I => \N__35137\
        );

    \I__6870\ : Span4Mux_h
    port map (
            O => \N__35137\,
            I => \N__35134\
        );

    \I__6869\ : Odrv4
    port map (
            O => \N__35134\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12\
        );

    \I__6868\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35127\
        );

    \I__6867\ : CascadeMux
    port map (
            O => \N__35130\,
            I => \N__35124\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__35127\,
            I => \N__35120\
        );

    \I__6865\ : InMux
    port map (
            O => \N__35124\,
            I => \N__35117\
        );

    \I__6864\ : InMux
    port map (
            O => \N__35123\,
            I => \N__35114\
        );

    \I__6863\ : Span4Mux_v
    port map (
            O => \N__35120\,
            I => \N__35111\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__35117\,
            I => \N__35108\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__35114\,
            I => \N__35105\
        );

    \I__6860\ : Span4Mux_h
    port map (
            O => \N__35111\,
            I => \N__35098\
        );

    \I__6859\ : Span4Mux_h
    port map (
            O => \N__35108\,
            I => \N__35098\
        );

    \I__6858\ : Span4Mux_h
    port map (
            O => \N__35105\,
            I => \N__35095\
        );

    \I__6857\ : InMux
    port map (
            O => \N__35104\,
            I => \N__35092\
        );

    \I__6856\ : InMux
    port map (
            O => \N__35103\,
            I => \N__35089\
        );

    \I__6855\ : Odrv4
    port map (
            O => \N__35098\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__6854\ : Odrv4
    port map (
            O => \N__35095\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__35092\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__35089\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__6851\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35075\
        );

    \I__6850\ : InMux
    port map (
            O => \N__35079\,
            I => \N__35072\
        );

    \I__6849\ : InMux
    port map (
            O => \N__35078\,
            I => \N__35069\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__35075\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__35072\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__35069\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\
        );

    \I__6845\ : InMux
    port map (
            O => \N__35062\,
            I => \N__35059\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__35059\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\
        );

    \I__6843\ : CascadeMux
    port map (
            O => \N__35056\,
            I => \N__35053\
        );

    \I__6842\ : InMux
    port map (
            O => \N__35053\,
            I => \N__35050\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__35050\,
            I => \N__35047\
        );

    \I__6840\ : Span4Mux_h
    port map (
            O => \N__35047\,
            I => \N__35044\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__35044\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0\
        );

    \I__6838\ : InMux
    port map (
            O => \N__35041\,
            I => \N__35037\
        );

    \I__6837\ : InMux
    port map (
            O => \N__35040\,
            I => \N__35033\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__35037\,
            I => \N__35030\
        );

    \I__6835\ : InMux
    port map (
            O => \N__35036\,
            I => \N__35027\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__35033\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__35030\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__35027\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\
        );

    \I__6831\ : InMux
    port map (
            O => \N__35020\,
            I => \N__35015\
        );

    \I__6830\ : InMux
    port map (
            O => \N__35019\,
            I => \N__35012\
        );

    \I__6829\ : InMux
    port map (
            O => \N__35018\,
            I => \N__35009\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__35015\,
            I => \N__35004\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__35012\,
            I => \N__35004\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__35009\,
            I => \N__35001\
        );

    \I__6825\ : Span4Mux_h
    port map (
            O => \N__35004\,
            I => \N__34998\
        );

    \I__6824\ : Odrv12
    port map (
            O => \N__35001\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6823\ : Odrv4
    port map (
            O => \N__34998\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6822\ : InMux
    port map (
            O => \N__34993\,
            I => \N__34990\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__34990\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\
        );

    \I__6820\ : InMux
    port map (
            O => \N__34987\,
            I => \N__34984\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__34984\,
            I => \N__34980\
        );

    \I__6818\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34976\
        );

    \I__6817\ : Span4Mux_h
    port map (
            O => \N__34980\,
            I => \N__34973\
        );

    \I__6816\ : InMux
    port map (
            O => \N__34979\,
            I => \N__34970\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__34976\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__34973\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__34970\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\
        );

    \I__6812\ : CascadeMux
    port map (
            O => \N__34963\,
            I => \N__34958\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34950\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34961\,
            I => \N__34950\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34950\
        );

    \I__6808\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34947\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__34950\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__34947\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6805\ : IoInMux
    port map (
            O => \N__34942\,
            I => \N__34939\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__34939\,
            I => \N__34936\
        );

    \I__6803\ : Span12Mux_s6_v
    port map (
            O => \N__34936\,
            I => \N__34931\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34926\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34934\,
            I => \N__34926\
        );

    \I__6800\ : Odrv12
    port map (
            O => \N__34931\,
            I => s1_phy_c
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__34926\,
            I => s1_phy_c
        );

    \I__6798\ : InMux
    port map (
            O => \N__34921\,
            I => \N__34915\
        );

    \I__6797\ : InMux
    port map (
            O => \N__34920\,
            I => \N__34910\
        );

    \I__6796\ : InMux
    port map (
            O => \N__34919\,
            I => \N__34910\
        );

    \I__6795\ : InMux
    port map (
            O => \N__34918\,
            I => \N__34907\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34915\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__34910\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__34907\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6791\ : IoInMux
    port map (
            O => \N__34900\,
            I => \N__34897\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__34897\,
            I => \N__34894\
        );

    \I__6789\ : Span4Mux_s3_v
    port map (
            O => \N__34894\,
            I => \N__34891\
        );

    \I__6788\ : Span4Mux_h
    port map (
            O => \N__34891\,
            I => \N__34887\
        );

    \I__6787\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34884\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__34887\,
            I => \T23_c\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__34884\,
            I => \T23_c\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34879\,
            I => \N__34874\
        );

    \I__6783\ : InMux
    port map (
            O => \N__34878\,
            I => \N__34870\
        );

    \I__6782\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34867\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34874\,
            I => \N__34864\
        );

    \I__6780\ : InMux
    port map (
            O => \N__34873\,
            I => \N__34861\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__34870\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__34867\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6777\ : Odrv12
    port map (
            O => \N__34864\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__34861\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6775\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34844\
        );

    \I__6774\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34844\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34841\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34838\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__34844\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__34841\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__34838\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6768\ : IoInMux
    port map (
            O => \N__34831\,
            I => \N__34828\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__34828\,
            I => \N__34825\
        );

    \I__6766\ : Odrv12
    port map (
            O => \N__34825\,
            I => \current_shift_inst.timer_s1.N_166_i\
        );

    \I__6765\ : IoInMux
    port map (
            O => \N__34822\,
            I => \N__34819\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__34819\,
            I => \N__34816\
        );

    \I__6763\ : Odrv12
    port map (
            O => \N__34816\,
            I => s2_phy_c
        );

    \I__6762\ : InMux
    port map (
            O => \N__34813\,
            I => \N__34810\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__34810\,
            I => \N__34807\
        );

    \I__6760\ : Span4Mux_h
    port map (
            O => \N__34807\,
            I => \N__34804\
        );

    \I__6759\ : Odrv4
    port map (
            O => \N__34804\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__34801\,
            I => \N__34798\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34793\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34790\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34796\,
            I => \N__34787\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__34793\,
            I => \N__34784\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__34790\,
            I => \N__34779\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__34787\,
            I => \N__34779\
        );

    \I__6751\ : Span4Mux_v
    port map (
            O => \N__34784\,
            I => \N__34776\
        );

    \I__6750\ : Span4Mux_v
    port map (
            O => \N__34779\,
            I => \N__34771\
        );

    \I__6749\ : Span4Mux_v
    port map (
            O => \N__34776\,
            I => \N__34768\
        );

    \I__6748\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34763\
        );

    \I__6747\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34763\
        );

    \I__6746\ : Sp12to4
    port map (
            O => \N__34771\,
            I => \N__34756\
        );

    \I__6745\ : Sp12to4
    port map (
            O => \N__34768\,
            I => \N__34756\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__34763\,
            I => \N__34756\
        );

    \I__6743\ : Odrv12
    port map (
            O => \N__34756\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34753\,
            I => \N__34750\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__34750\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\
        );

    \I__6740\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34743\
        );

    \I__6739\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34740\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__34743\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__34740\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\
        );

    \I__6736\ : InMux
    port map (
            O => \N__34735\,
            I => \N__34731\
        );

    \I__6735\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34728\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__34731\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__34728\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\
        );

    \I__6732\ : CascadeMux
    port map (
            O => \N__34723\,
            I => \elapsed_time_ns_1_RNIP93CP1_0_1_cascade_\
        );

    \I__6731\ : CascadeMux
    port map (
            O => \N__34720\,
            I => \N__34716\
        );

    \I__6730\ : InMux
    port map (
            O => \N__34719\,
            I => \N__34713\
        );

    \I__6729\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34710\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__34713\,
            I => \N__34705\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__34710\,
            I => \N__34705\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__34705\,
            I => \phase_controller_inst1.stoper_hc.N_310\
        );

    \I__6725\ : CascadeMux
    port map (
            O => \N__34702\,
            I => \N__34698\
        );

    \I__6724\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34695\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34692\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__34695\,
            I => \N__34689\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__34692\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__34689\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\
        );

    \I__6719\ : CascadeMux
    port map (
            O => \N__34684\,
            I => \N__34681\
        );

    \I__6718\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34678\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__34678\,
            I => \N__34675\
        );

    \I__6716\ : Odrv4
    port map (
            O => \N__34675\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__6715\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34668\
        );

    \I__6714\ : InMux
    port map (
            O => \N__34671\,
            I => \N__34665\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__34668\,
            I => state_ns_i_a2_1
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__34665\,
            I => state_ns_i_a2_1
        );

    \I__6711\ : InMux
    port map (
            O => \N__34660\,
            I => \N__34656\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34653\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__34656\,
            I => \N__34650\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__34653\,
            I => \N__34646\
        );

    \I__6707\ : Span4Mux_v
    port map (
            O => \N__34650\,
            I => \N__34643\
        );

    \I__6706\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34640\
        );

    \I__6705\ : Span12Mux_s9_v
    port map (
            O => \N__34646\,
            I => \N__34637\
        );

    \I__6704\ : Odrv4
    port map (
            O => \N__34643\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__34640\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6702\ : Odrv12
    port map (
            O => \N__34637\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6701\ : IoInMux
    port map (
            O => \N__34630\,
            I => \N__34627\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__34627\,
            I => \N__34624\
        );

    \I__6699\ : Span4Mux_s3_v
    port map (
            O => \N__34624\,
            I => \N__34621\
        );

    \I__6698\ : Span4Mux_v
    port map (
            O => \N__34621\,
            I => \N__34617\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34620\,
            I => \N__34614\
        );

    \I__6696\ : Odrv4
    port map (
            O => \N__34617\,
            I => \T45_c\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__34614\,
            I => \T45_c\
        );

    \I__6694\ : CascadeMux
    port map (
            O => \N__34609\,
            I => \N__34604\
        );

    \I__6693\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34601\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__34607\,
            I => \N__34598\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34604\,
            I => \N__34594\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__34601\,
            I => \N__34591\
        );

    \I__6689\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34588\
        );

    \I__6688\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34585\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__34594\,
            I => \elapsed_time_ns_1_RNIRB3CP1_0_3\
        );

    \I__6686\ : Odrv4
    port map (
            O => \N__34591\,
            I => \elapsed_time_ns_1_RNIRB3CP1_0_3\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__34588\,
            I => \elapsed_time_ns_1_RNIRB3CP1_0_3\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__34585\,
            I => \elapsed_time_ns_1_RNIRB3CP1_0_3\
        );

    \I__6683\ : CascadeMux
    port map (
            O => \N__34576\,
            I => \N__34573\
        );

    \I__6682\ : InMux
    port map (
            O => \N__34573\,
            I => \N__34564\
        );

    \I__6681\ : InMux
    port map (
            O => \N__34572\,
            I => \N__34564\
        );

    \I__6680\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34564\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__34564\,
            I => \elapsed_time_ns_1_RNIJEKEE1_0_2\
        );

    \I__6678\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34558\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__34558\,
            I => \phase_controller_inst1.stoper_hc.N_286\
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__34555\,
            I => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1_cascade_\
        );

    \I__6675\ : InMux
    port map (
            O => \N__34552\,
            I => \N__34546\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34551\,
            I => \N__34546\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__34546\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__6672\ : CascadeMux
    port map (
            O => \N__34543\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_\
        );

    \I__6671\ : CascadeMux
    port map (
            O => \N__34540\,
            I => \phase_controller_inst1.stoper_hc.N_328_cascade_\
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__34537\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\
        );

    \I__6669\ : InMux
    port map (
            O => \N__34534\,
            I => \N__34529\
        );

    \I__6668\ : InMux
    port map (
            O => \N__34533\,
            I => \N__34524\
        );

    \I__6667\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34524\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__34529\,
            I => \elapsed_time_ns_1_RNIP93CP1_0_1\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__34524\,
            I => \elapsed_time_ns_1_RNIP93CP1_0_1\
        );

    \I__6664\ : InMux
    port map (
            O => \N__34519\,
            I => \N__34515\
        );

    \I__6663\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34512\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__34515\,
            I => \N__34507\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__34512\,
            I => \N__34507\
        );

    \I__6660\ : Span4Mux_v
    port map (
            O => \N__34507\,
            I => \N__34502\
        );

    \I__6659\ : InMux
    port map (
            O => \N__34506\,
            I => \N__34497\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34505\,
            I => \N__34497\
        );

    \I__6657\ : Odrv4
    port map (
            O => \N__34502\,
            I => \elapsed_time_ns_1_RNIPKKEE1_0_8\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__34497\,
            I => \elapsed_time_ns_1_RNIPKKEE1_0_8\
        );

    \I__6655\ : CascadeMux
    port map (
            O => \N__34492\,
            I => \elapsed_time_ns_1_RNIOJKEE1_0_7_cascade_\
        );

    \I__6654\ : CascadeMux
    port map (
            O => \N__34489\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\
        );

    \I__6653\ : CascadeMux
    port map (
            O => \N__34486\,
            I => \phase_controller_inst1.stoper_hc.N_330_cascade_\
        );

    \I__6652\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34479\
        );

    \I__6651\ : InMux
    port map (
            O => \N__34482\,
            I => \N__34476\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__34479\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__34476\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\
        );

    \I__6648\ : InMux
    port map (
            O => \N__34471\,
            I => \N__34467\
        );

    \I__6647\ : InMux
    port map (
            O => \N__34470\,
            I => \N__34464\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__34467\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__34464\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2\
        );

    \I__6644\ : CascadeMux
    port map (
            O => \N__34459\,
            I => \N__34456\
        );

    \I__6643\ : InMux
    port map (
            O => \N__34456\,
            I => \N__34451\
        );

    \I__6642\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34446\
        );

    \I__6641\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34446\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__34451\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__34446\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\
        );

    \I__6638\ : CascadeMux
    port map (
            O => \N__34441\,
            I => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34438\,
            I => \N__34435\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__34435\,
            I => \N__34432\
        );

    \I__6635\ : Odrv12
    port map (
            O => \N__34432\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df28\
        );

    \I__6634\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34426\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__34426\,
            I => \N__34423\
        );

    \I__6632\ : Odrv12
    port map (
            O => \N__34423\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__6631\ : InMux
    port map (
            O => \N__34420\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28\
        );

    \I__6630\ : InMux
    port map (
            O => \N__34417\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__6629\ : CascadeMux
    port map (
            O => \N__34414\,
            I => \N__34411\
        );

    \I__6628\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34408\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__34408\,
            I => \N__34405\
        );

    \I__6626\ : Odrv12
    port map (
            O => \N__34405\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__6625\ : InMux
    port map (
            O => \N__34402\,
            I => \N__34399\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__34399\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__6623\ : InMux
    port map (
            O => \N__34396\,
            I => \N__34393\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__34393\,
            I => \N__34390\
        );

    \I__6621\ : Odrv12
    port map (
            O => \N__34390\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__6620\ : CascadeMux
    port map (
            O => \N__34387\,
            I => \N__34384\
        );

    \I__6619\ : InMux
    port map (
            O => \N__34384\,
            I => \N__34381\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__34381\,
            I => \N__34378\
        );

    \I__6617\ : Odrv4
    port map (
            O => \N__34378\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__6616\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34372\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__34372\,
            I => \N__34369\
        );

    \I__6614\ : Odrv12
    port map (
            O => \N__34369\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__6613\ : CascadeMux
    port map (
            O => \N__34366\,
            I => \N__34363\
        );

    \I__6612\ : InMux
    port map (
            O => \N__34363\,
            I => \N__34360\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__34360\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__6610\ : InMux
    port map (
            O => \N__34357\,
            I => \N__34354\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__34354\,
            I => \N__34351\
        );

    \I__6608\ : Odrv12
    port map (
            O => \N__34351\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__6607\ : CascadeMux
    port map (
            O => \N__34348\,
            I => \N__34345\
        );

    \I__6606\ : InMux
    port map (
            O => \N__34345\,
            I => \N__34342\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__34342\,
            I => \N__34339\
        );

    \I__6604\ : Odrv4
    port map (
            O => \N__34339\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__6603\ : InMux
    port map (
            O => \N__34336\,
            I => \N__34333\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__34333\,
            I => \N__34330\
        );

    \I__6601\ : Odrv12
    port map (
            O => \N__34330\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__6600\ : CascadeMux
    port map (
            O => \N__34327\,
            I => \N__34324\
        );

    \I__6599\ : InMux
    port map (
            O => \N__34324\,
            I => \N__34321\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__34321\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__6597\ : CascadeMux
    port map (
            O => \N__34318\,
            I => \N__34315\
        );

    \I__6596\ : InMux
    port map (
            O => \N__34315\,
            I => \N__34312\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__34312\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__6594\ : CascadeMux
    port map (
            O => \N__34309\,
            I => \N__34306\
        );

    \I__6593\ : InMux
    port map (
            O => \N__34306\,
            I => \N__34303\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__34303\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__6591\ : InMux
    port map (
            O => \N__34300\,
            I => \N__34297\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__34297\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__6589\ : CascadeMux
    port map (
            O => \N__34294\,
            I => \N__34291\
        );

    \I__6588\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34288\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__34288\,
            I => \N__34285\
        );

    \I__6586\ : Odrv4
    port map (
            O => \N__34285\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__6585\ : InMux
    port map (
            O => \N__34282\,
            I => \N__34279\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__34279\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__6583\ : CascadeMux
    port map (
            O => \N__34276\,
            I => \N__34273\
        );

    \I__6582\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34270\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__34270\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__6580\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34264\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__34264\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__6578\ : CascadeMux
    port map (
            O => \N__34261\,
            I => \N__34258\
        );

    \I__6577\ : InMux
    port map (
            O => \N__34258\,
            I => \N__34255\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__34255\,
            I => \N__34252\
        );

    \I__6575\ : Odrv4
    port map (
            O => \N__34252\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__6574\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34246\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__34246\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__6572\ : CascadeMux
    port map (
            O => \N__34243\,
            I => \N__34240\
        );

    \I__6571\ : InMux
    port map (
            O => \N__34240\,
            I => \N__34237\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__34237\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__6569\ : CascadeMux
    port map (
            O => \N__34234\,
            I => \N__34231\
        );

    \I__6568\ : InMux
    port map (
            O => \N__34231\,
            I => \N__34228\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__34228\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__6566\ : InMux
    port map (
            O => \N__34225\,
            I => \N__34222\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__34222\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__6564\ : CascadeMux
    port map (
            O => \N__34219\,
            I => \N__34216\
        );

    \I__6563\ : InMux
    port map (
            O => \N__34216\,
            I => \N__34213\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__34213\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__6561\ : InMux
    port map (
            O => \N__34210\,
            I => \N__34207\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__34207\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__6559\ : InMux
    port map (
            O => \N__34204\,
            I => \N__34201\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__34201\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__6557\ : IoInMux
    port map (
            O => \N__34198\,
            I => \N__34195\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__34195\,
            I => \N__34192\
        );

    \I__6555\ : IoSpan4Mux
    port map (
            O => \N__34192\,
            I => \N__34189\
        );

    \I__6554\ : Span4Mux_s1_v
    port map (
            O => \N__34189\,
            I => \N__34186\
        );

    \I__6553\ : Sp12to4
    port map (
            O => \N__34186\,
            I => \N__34183\
        );

    \I__6552\ : Span12Mux_s9_v
    port map (
            O => \N__34183\,
            I => \N__34180\
        );

    \I__6551\ : Odrv12
    port map (
            O => \N__34180\,
            I => \pll_inst.red_c_i\
        );

    \I__6550\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34174\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__34174\,
            I => \N__34169\
        );

    \I__6548\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34166\
        );

    \I__6547\ : InMux
    port map (
            O => \N__34172\,
            I => \N__34163\
        );

    \I__6546\ : Sp12to4
    port map (
            O => \N__34169\,
            I => \N__34158\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__34166\,
            I => \N__34158\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__34163\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__6543\ : Odrv12
    port map (
            O => \N__34158\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\
        );

    \I__6542\ : CascadeMux
    port map (
            O => \N__34153\,
            I => \N__34150\
        );

    \I__6541\ : InMux
    port map (
            O => \N__34150\,
            I => \N__34147\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__34147\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__6539\ : InMux
    port map (
            O => \N__34144\,
            I => \N__34141\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__34141\,
            I => \N__34136\
        );

    \I__6537\ : InMux
    port map (
            O => \N__34140\,
            I => \N__34133\
        );

    \I__6536\ : InMux
    port map (
            O => \N__34139\,
            I => \N__34130\
        );

    \I__6535\ : Sp12to4
    port map (
            O => \N__34136\,
            I => \N__34125\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__34133\,
            I => \N__34125\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__34130\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__6532\ : Odrv12
    port map (
            O => \N__34125\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\
        );

    \I__6531\ : InMux
    port map (
            O => \N__34120\,
            I => \N__34117\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__34117\,
            I => \N__34114\
        );

    \I__6529\ : Odrv4
    port map (
            O => \N__34114\,
            I => \current_shift_inst.PI_CTRL.integrator_i_24\
        );

    \I__6528\ : InMux
    port map (
            O => \N__34111\,
            I => \N__34106\
        );

    \I__6527\ : InMux
    port map (
            O => \N__34110\,
            I => \N__34103\
        );

    \I__6526\ : InMux
    port map (
            O => \N__34109\,
            I => \N__34100\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__34106\,
            I => \N__34097\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__34103\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__34100\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__6522\ : Odrv12
    port map (
            O => \N__34097\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__34090\,
            I => \N__34087\
        );

    \I__6520\ : InMux
    port map (
            O => \N__34087\,
            I => \N__34081\
        );

    \I__6519\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34078\
        );

    \I__6518\ : InMux
    port map (
            O => \N__34085\,
            I => \N__34075\
        );

    \I__6517\ : InMux
    port map (
            O => \N__34084\,
            I => \N__34072\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__34081\,
            I => \N__34069\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__34078\,
            I => \N__34066\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__34075\,
            I => \N__34061\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__34072\,
            I => \N__34061\
        );

    \I__6512\ : Span4Mux_h
    port map (
            O => \N__34069\,
            I => \N__34057\
        );

    \I__6511\ : Span4Mux_v
    port map (
            O => \N__34066\,
            I => \N__34052\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__34061\,
            I => \N__34052\
        );

    \I__6509\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34049\
        );

    \I__6508\ : Odrv4
    port map (
            O => \N__34057\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__6507\ : Odrv4
    port map (
            O => \N__34052\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__34049\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__6505\ : InMux
    port map (
            O => \N__34042\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_31\
        );

    \I__6504\ : InMux
    port map (
            O => \N__34039\,
            I => \N__34036\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__34036\,
            I => \N__34033\
        );

    \I__6502\ : Span4Mux_h
    port map (
            O => \N__34033\,
            I => \N__34030\
        );

    \I__6501\ : Odrv4
    port map (
            O => \N__34030\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0\
        );

    \I__6500\ : CascadeMux
    port map (
            O => \N__34027\,
            I => \N__34024\
        );

    \I__6499\ : InMux
    port map (
            O => \N__34024\,
            I => \N__34021\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__34021\,
            I => \N__34018\
        );

    \I__6497\ : Odrv12
    port map (
            O => \N__34018\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__6496\ : CascadeMux
    port map (
            O => \N__34015\,
            I => \N__34012\
        );

    \I__6495\ : InMux
    port map (
            O => \N__34012\,
            I => \N__34008\
        );

    \I__6494\ : CascadeMux
    port map (
            O => \N__34011\,
            I => \N__34003\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__34008\,
            I => \N__33999\
        );

    \I__6492\ : InMux
    port map (
            O => \N__34007\,
            I => \N__33994\
        );

    \I__6491\ : InMux
    port map (
            O => \N__34006\,
            I => \N__33994\
        );

    \I__6490\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33989\
        );

    \I__6489\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33989\
        );

    \I__6488\ : Span12Mux_v
    port map (
            O => \N__33999\,
            I => \N__33984\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__33994\,
            I => \N__33984\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33989\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__6485\ : Odrv12
    port map (
            O => \N__33984\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__6484\ : CascadeMux
    port map (
            O => \N__33979\,
            I => \N__33976\
        );

    \I__6483\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33973\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__33973\,
            I => \N__33970\
        );

    \I__6481\ : Odrv4
    port map (
            O => \N__33970\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33967\,
            I => \N__33964\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__33964\,
            I => \N__33961\
        );

    \I__6478\ : Span4Mux_h
    port map (
            O => \N__33961\,
            I => \N__33958\
        );

    \I__6477\ : Odrv4
    port map (
            O => \N__33958\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__6476\ : CascadeMux
    port map (
            O => \N__33955\,
            I => \N__33952\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33952\,
            I => \N__33946\
        );

    \I__6474\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33943\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33940\
        );

    \I__6472\ : InMux
    port map (
            O => \N__33949\,
            I => \N__33937\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33946\,
            I => \N__33933\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__33943\,
            I => \N__33930\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__33940\,
            I => \N__33927\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__33937\,
            I => \N__33924\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33921\
        );

    \I__6466\ : Span4Mux_v
    port map (
            O => \N__33933\,
            I => \N__33918\
        );

    \I__6465\ : Span4Mux_v
    port map (
            O => \N__33930\,
            I => \N__33911\
        );

    \I__6464\ : Span4Mux_v
    port map (
            O => \N__33927\,
            I => \N__33911\
        );

    \I__6463\ : Span4Mux_v
    port map (
            O => \N__33924\,
            I => \N__33911\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__33921\,
            I => \N__33908\
        );

    \I__6461\ : Span4Mux_h
    port map (
            O => \N__33918\,
            I => \N__33905\
        );

    \I__6460\ : Span4Mux_h
    port map (
            O => \N__33911\,
            I => \N__33902\
        );

    \I__6459\ : Odrv12
    port map (
            O => \N__33908\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__6458\ : Odrv4
    port map (
            O => \N__33905\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__6457\ : Odrv4
    port map (
            O => \N__33902\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__6456\ : CascadeMux
    port map (
            O => \N__33895\,
            I => \N__33892\
        );

    \I__6455\ : InMux
    port map (
            O => \N__33892\,
            I => \N__33889\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__33889\,
            I => \N__33886\
        );

    \I__6453\ : Odrv4
    port map (
            O => \N__33886\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__6452\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33880\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__33880\,
            I => \N__33877\
        );

    \I__6450\ : Span4Mux_h
    port map (
            O => \N__33877\,
            I => \N__33874\
        );

    \I__6449\ : Odrv4
    port map (
            O => \N__33874\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__33871\,
            I => \N__33868\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33868\,
            I => \N__33864\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33867\,
            I => \N__33859\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__33864\,
            I => \N__33856\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33853\
        );

    \I__6443\ : InMux
    port map (
            O => \N__33862\,
            I => \N__33850\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__33859\,
            I => \N__33847\
        );

    \I__6441\ : Span4Mux_v
    port map (
            O => \N__33856\,
            I => \N__33844\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__33853\,
            I => \N__33841\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__33850\,
            I => \N__33837\
        );

    \I__6438\ : Span4Mux_v
    port map (
            O => \N__33847\,
            I => \N__33832\
        );

    \I__6437\ : Span4Mux_h
    port map (
            O => \N__33844\,
            I => \N__33832\
        );

    \I__6436\ : Span4Mux_v
    port map (
            O => \N__33841\,
            I => \N__33829\
        );

    \I__6435\ : InMux
    port map (
            O => \N__33840\,
            I => \N__33826\
        );

    \I__6434\ : Odrv12
    port map (
            O => \N__33837\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__6433\ : Odrv4
    port map (
            O => \N__33832\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__6432\ : Odrv4
    port map (
            O => \N__33829\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__33826\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__6430\ : InMux
    port map (
            O => \N__33817\,
            I => \N__33814\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__33814\,
            I => \N__33809\
        );

    \I__6428\ : CascadeMux
    port map (
            O => \N__33813\,
            I => \N__33806\
        );

    \I__6427\ : CascadeMux
    port map (
            O => \N__33812\,
            I => \N__33803\
        );

    \I__6426\ : Span4Mux_h
    port map (
            O => \N__33809\,
            I => \N__33799\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33806\,
            I => \N__33796\
        );

    \I__6424\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33793\
        );

    \I__6423\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33789\
        );

    \I__6422\ : Span4Mux_h
    port map (
            O => \N__33799\,
            I => \N__33786\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__33796\,
            I => \N__33781\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__33793\,
            I => \N__33781\
        );

    \I__6419\ : InMux
    port map (
            O => \N__33792\,
            I => \N__33778\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__33789\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6417\ : Odrv4
    port map (
            O => \N__33786\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6416\ : Odrv12
    port map (
            O => \N__33781\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__33778\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__33769\,
            I => \N__33766\
        );

    \I__6413\ : InMux
    port map (
            O => \N__33766\,
            I => \N__33763\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__33763\,
            I => \N__33760\
        );

    \I__6411\ : Span4Mux_v
    port map (
            O => \N__33760\,
            I => \N__33757\
        );

    \I__6410\ : Odrv4
    port map (
            O => \N__33757\,
            I => \current_shift_inst.PI_CTRL.integrator_i_21\
        );

    \I__6409\ : CascadeMux
    port map (
            O => \N__33754\,
            I => \N__33750\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33753\,
            I => \N__33747\
        );

    \I__6407\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33744\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__33747\,
            I => \N__33740\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__33744\,
            I => \N__33737\
        );

    \I__6404\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33734\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__33740\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__6402\ : Odrv12
    port map (
            O => \N__33737\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__33734\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__6400\ : InMux
    port map (
            O => \N__33727\,
            I => \N__33724\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__33724\,
            I => \N__33721\
        );

    \I__6398\ : Odrv12
    port map (
            O => \N__33721\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\
        );

    \I__6397\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33713\
        );

    \I__6396\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33710\
        );

    \I__6395\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33707\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__33713\,
            I => \N__33704\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__33710\,
            I => \N__33699\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33707\,
            I => \N__33696\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__33704\,
            I => \N__33693\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33688\
        );

    \I__6389\ : InMux
    port map (
            O => \N__33702\,
            I => \N__33688\
        );

    \I__6388\ : Span4Mux_h
    port map (
            O => \N__33699\,
            I => \N__33685\
        );

    \I__6387\ : Odrv4
    port map (
            O => \N__33696\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__6386\ : Odrv4
    port map (
            O => \N__33693\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__33688\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__6384\ : Odrv4
    port map (
            O => \N__33685\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33673\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__33673\,
            I => \N__33670\
        );

    \I__6381\ : Span4Mux_h
    port map (
            O => \N__33670\,
            I => \N__33667\
        );

    \I__6380\ : Odrv4
    port map (
            O => \N__33667\,
            I => \current_shift_inst.PI_CTRL.integrator_i_17\
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__33664\,
            I => \N__33661\
        );

    \I__6378\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33658\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__33658\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\
        );

    \I__6376\ : InMux
    port map (
            O => \N__33655\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\
        );

    \I__6375\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33649\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__33649\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\
        );

    \I__6373\ : InMux
    port map (
            O => \N__33646\,
            I => \bfn_13_7_0_\
        );

    \I__6372\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33639\
        );

    \I__6371\ : InMux
    port map (
            O => \N__33642\,
            I => \N__33636\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__33639\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__33636\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\
        );

    \I__6368\ : InMux
    port map (
            O => \N__33631\,
            I => \N__33628\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__33628\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\
        );

    \I__6366\ : InMux
    port map (
            O => \N__33625\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\
        );

    \I__6365\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33619\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__33619\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\
        );

    \I__6363\ : InMux
    port map (
            O => \N__33616\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\
        );

    \I__6362\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33610\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__33610\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\
        );

    \I__6360\ : InMux
    port map (
            O => \N__33607\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\
        );

    \I__6359\ : InMux
    port map (
            O => \N__33604\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\
        );

    \I__6358\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33598\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__33598\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\
        );

    \I__6356\ : InMux
    port map (
            O => \N__33595\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\
        );

    \I__6355\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33589\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__33589\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\
        );

    \I__6353\ : InMux
    port map (
            O => \N__33586\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__33583\,
            I => \N__33580\
        );

    \I__6351\ : InMux
    port map (
            O => \N__33580\,
            I => \N__33577\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__33577\,
            I => \N__33574\
        );

    \I__6349\ : Odrv4
    port map (
            O => \N__33574\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\
        );

    \I__6348\ : InMux
    port map (
            O => \N__33571\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\
        );

    \I__6347\ : InMux
    port map (
            O => \N__33568\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\
        );

    \I__6346\ : InMux
    port map (
            O => \N__33565\,
            I => \N__33562\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__33562\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\
        );

    \I__6344\ : InMux
    port map (
            O => \N__33559\,
            I => \bfn_13_6_0_\
        );

    \I__6343\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33553\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__33553\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\
        );

    \I__6341\ : InMux
    port map (
            O => \N__33550\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33542\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33546\,
            I => \N__33539\
        );

    \I__6338\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33536\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__33542\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__33539\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__33536\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\
        );

    \I__6334\ : CascadeMux
    port map (
            O => \N__33529\,
            I => \N__33526\
        );

    \I__6333\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33523\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33520\
        );

    \I__6331\ : Odrv4
    port map (
            O => \N__33520\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\
        );

    \I__6330\ : InMux
    port map (
            O => \N__33517\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__33514\,
            I => \N__33511\
        );

    \I__6328\ : InMux
    port map (
            O => \N__33511\,
            I => \N__33508\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__33508\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\
        );

    \I__6326\ : InMux
    port map (
            O => \N__33505\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\
        );

    \I__6325\ : InMux
    port map (
            O => \N__33502\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\
        );

    \I__6324\ : InMux
    port map (
            O => \N__33499\,
            I => \N__33496\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__33496\,
            I => \N__33493\
        );

    \I__6322\ : Odrv4
    port map (
            O => \N__33493\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\
        );

    \I__6321\ : InMux
    port map (
            O => \N__33490\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\
        );

    \I__6320\ : InMux
    port map (
            O => \N__33487\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\
        );

    \I__6319\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33481\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__33481\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\
        );

    \I__6317\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33475\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__33475\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_6\
        );

    \I__6315\ : InMux
    port map (
            O => \N__33472\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\
        );

    \I__6314\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33466\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__33466\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\
        );

    \I__6312\ : CascadeMux
    port map (
            O => \N__33463\,
            I => \N__33460\
        );

    \I__6311\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33457\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__33457\,
            I => \N__33454\
        );

    \I__6309\ : Odrv4
    port map (
            O => \N__33454\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_7\
        );

    \I__6308\ : InMux
    port map (
            O => \N__33451\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\
        );

    \I__6307\ : InMux
    port map (
            O => \N__33448\,
            I => \N__33445\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__33445\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\
        );

    \I__6305\ : InMux
    port map (
            O => \N__33442\,
            I => \N__33439\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__33439\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_8\
        );

    \I__6303\ : InMux
    port map (
            O => \N__33436\,
            I => \bfn_13_5_0_\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__33433\,
            I => \N__33430\
        );

    \I__6301\ : InMux
    port map (
            O => \N__33430\,
            I => \N__33427\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__33427\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_9\
        );

    \I__6299\ : InMux
    port map (
            O => \N__33424\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\
        );

    \I__6298\ : InMux
    port map (
            O => \N__33421\,
            I => \N__33418\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__33418\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\
        );

    \I__6296\ : CascadeMux
    port map (
            O => \N__33415\,
            I => \N__33412\
        );

    \I__6295\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33409\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__33409\,
            I => \N__33406\
        );

    \I__6293\ : Odrv4
    port map (
            O => \N__33406\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_10\
        );

    \I__6292\ : InMux
    port map (
            O => \N__33403\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\
        );

    \I__6291\ : InMux
    port map (
            O => \N__33400\,
            I => \N__33397\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__33397\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\
        );

    \I__6289\ : CascadeMux
    port map (
            O => \N__33394\,
            I => \N__33391\
        );

    \I__6288\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33388\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__33388\,
            I => \N__33385\
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__33385\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_11\
        );

    \I__6285\ : InMux
    port map (
            O => \N__33382\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\
        );

    \I__6284\ : InMux
    port map (
            O => \N__33379\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\
        );

    \I__6283\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33373\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__33373\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_13\
        );

    \I__6281\ : InMux
    port map (
            O => \N__33370\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\
        );

    \I__6280\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33361\
        );

    \I__6279\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33361\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__33361\,
            I => \phase_controller_inst1.N_54\
        );

    \I__6277\ : CEMux
    port map (
            O => \N__33358\,
            I => \N__33353\
        );

    \I__6276\ : CEMux
    port map (
            O => \N__33357\,
            I => \N__33350\
        );

    \I__6275\ : CEMux
    port map (
            O => \N__33356\,
            I => \N__33347\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__33353\,
            I => \N__33342\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__33350\,
            I => \N__33342\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__33347\,
            I => \N__33338\
        );

    \I__6271\ : Span4Mux_v
    port map (
            O => \N__33342\,
            I => \N__33335\
        );

    \I__6270\ : CEMux
    port map (
            O => \N__33341\,
            I => \N__33332\
        );

    \I__6269\ : Span4Mux_v
    port map (
            O => \N__33338\,
            I => \N__33325\
        );

    \I__6268\ : Span4Mux_h
    port map (
            O => \N__33335\,
            I => \N__33325\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__33332\,
            I => \N__33325\
        );

    \I__6266\ : Span4Mux_h
    port map (
            O => \N__33325\,
            I => \N__33322\
        );

    \I__6265\ : Span4Mux_h
    port map (
            O => \N__33322\,
            I => \N__33319\
        );

    \I__6264\ : Odrv4
    port map (
            O => \N__33319\,
            I => \current_shift_inst.timer_s1.N_167_i\
        );

    \I__6263\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33313\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__33313\,
            I => \N__33309\
        );

    \I__6261\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33306\
        );

    \I__6260\ : Span4Mux_h
    port map (
            O => \N__33309\,
            I => \N__33303\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__33306\,
            I => \N__33298\
        );

    \I__6258\ : Span4Mux_v
    port map (
            O => \N__33303\,
            I => \N__33298\
        );

    \I__6257\ : Odrv4
    port map (
            O => \N__33298\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__6256\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33292\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__33292\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\
        );

    \I__6254\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33285\
        );

    \I__6253\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33282\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__33285\,
            I => \N__33279\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__33282\,
            I => \N__33276\
        );

    \I__6250\ : Span4Mux_v
    port map (
            O => \N__33279\,
            I => \N__33273\
        );

    \I__6249\ : Odrv4
    port map (
            O => \N__33276\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__6248\ : Odrv4
    port map (
            O => \N__33273\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__6247\ : CascadeMux
    port map (
            O => \N__33268\,
            I => \N__33265\
        );

    \I__6246\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33262\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__33262\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\
        );

    \I__6244\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33255\
        );

    \I__6243\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33252\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__33255\,
            I => \N__33249\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__33252\,
            I => \N__33246\
        );

    \I__6240\ : Span4Mux_v
    port map (
            O => \N__33249\,
            I => \N__33243\
        );

    \I__6239\ : Odrv4
    port map (
            O => \N__33246\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__6238\ : Odrv4
    port map (
            O => \N__33243\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__6237\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33235\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__33235\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\
        );

    \I__6235\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33228\
        );

    \I__6234\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33225\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__33228\,
            I => \N__33222\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__33225\,
            I => \N__33219\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__33222\,
            I => \N__33216\
        );

    \I__6230\ : Odrv12
    port map (
            O => \N__33219\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__33216\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6228\ : InMux
    port map (
            O => \N__33211\,
            I => \N__33208\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__33208\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\
        );

    \I__6226\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33202\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__33202\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\
        );

    \I__6224\ : InMux
    port map (
            O => \N__33199\,
            I => \N__33196\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__33196\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_4\
        );

    \I__6222\ : InMux
    port map (
            O => \N__33193\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\
        );

    \I__6221\ : InMux
    port map (
            O => \N__33190\,
            I => \N__33187\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__33187\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33181\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__33181\,
            I => \current_shift_inst.PI_CTRL.un7_integrator1_5\
        );

    \I__6217\ : InMux
    port map (
            O => \N__33178\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\
        );

    \I__6216\ : CascadeMux
    port map (
            O => \N__33175\,
            I => \N__33172\
        );

    \I__6215\ : InMux
    port map (
            O => \N__33172\,
            I => \N__33169\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__33169\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__6213\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33163\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__33163\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__6211\ : InMux
    port map (
            O => \N__33160\,
            I => \N__33157\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__33157\,
            I => \N__33153\
        );

    \I__6209\ : InMux
    port map (
            O => \N__33156\,
            I => \N__33150\
        );

    \I__6208\ : Span4Mux_s1_v
    port map (
            O => \N__33153\,
            I => \N__33144\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__33150\,
            I => \N__33144\
        );

    \I__6206\ : InMux
    port map (
            O => \N__33149\,
            I => \N__33141\
        );

    \I__6205\ : Span4Mux_v
    port map (
            O => \N__33144\,
            I => \N__33137\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__33141\,
            I => \N__33134\
        );

    \I__6203\ : InMux
    port map (
            O => \N__33140\,
            I => \N__33131\
        );

    \I__6202\ : Span4Mux_h
    port map (
            O => \N__33137\,
            I => \N__33128\
        );

    \I__6201\ : Span4Mux_v
    port map (
            O => \N__33134\,
            I => \N__33123\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__33131\,
            I => \N__33123\
        );

    \I__6199\ : Sp12to4
    port map (
            O => \N__33128\,
            I => \N__33120\
        );

    \I__6198\ : Span4Mux_v
    port map (
            O => \N__33123\,
            I => \N__33117\
        );

    \I__6197\ : Span12Mux_v
    port map (
            O => \N__33120\,
            I => \N__33114\
        );

    \I__6196\ : Span4Mux_v
    port map (
            O => \N__33117\,
            I => \N__33111\
        );

    \I__6195\ : Span12Mux_v
    port map (
            O => \N__33114\,
            I => \N__33108\
        );

    \I__6194\ : Sp12to4
    port map (
            O => \N__33111\,
            I => \N__33105\
        );

    \I__6193\ : Span12Mux_h
    port map (
            O => \N__33108\,
            I => \N__33102\
        );

    \I__6192\ : Span12Mux_h
    port map (
            O => \N__33105\,
            I => \N__33099\
        );

    \I__6191\ : Odrv12
    port map (
            O => \N__33102\,
            I => start_stop_c
        );

    \I__6190\ : Odrv12
    port map (
            O => \N__33099\,
            I => start_stop_c
        );

    \I__6189\ : InMux
    port map (
            O => \N__33094\,
            I => \N__33091\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__33091\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__6187\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33081\
        );

    \I__6186\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33072\
        );

    \I__6185\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33072\
        );

    \I__6184\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33072\
        );

    \I__6183\ : InMux
    port map (
            O => \N__33084\,
            I => \N__33072\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__33081\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__33072\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__33067\,
            I => \N__33063\
        );

    \I__6179\ : InMux
    port map (
            O => \N__33066\,
            I => \N__33056\
        );

    \I__6178\ : InMux
    port map (
            O => \N__33063\,
            I => \N__33056\
        );

    \I__6177\ : InMux
    port map (
            O => \N__33062\,
            I => \N__33053\
        );

    \I__6176\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33050\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__33056\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__33053\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__33050\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__6172\ : InMux
    port map (
            O => \N__33043\,
            I => \N__33040\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__33040\,
            I => \N__33037\
        );

    \I__6170\ : Span4Mux_v
    port map (
            O => \N__33037\,
            I => \N__33034\
        );

    \I__6169\ : Odrv4
    port map (
            O => \N__33034\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__6168\ : InMux
    port map (
            O => \N__33031\,
            I => \N__33028\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__33025\
        );

    \I__6166\ : Odrv4
    port map (
            O => \N__33025\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__6165\ : InMux
    port map (
            O => \N__33022\,
            I => \N__33019\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__33019\,
            I => \N__33016\
        );

    \I__6163\ : Sp12to4
    port map (
            O => \N__33016\,
            I => \N__33013\
        );

    \I__6162\ : Odrv12
    port map (
            O => \N__33013\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__6161\ : InMux
    port map (
            O => \N__33010\,
            I => \N__33007\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__33007\,
            I => \N__33004\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__33004\,
            I => \N__33001\
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__33001\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32998\,
            I => \N__32995\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__32995\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32992\,
            I => \N__32989\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__32989\,
            I => \N__32986\
        );

    \I__6153\ : Odrv12
    port map (
            O => \N__32986\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__6152\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32980\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__32980\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__6150\ : CascadeMux
    port map (
            O => \N__32977\,
            I => \N__32974\
        );

    \I__6149\ : InMux
    port map (
            O => \N__32974\,
            I => \N__32971\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__32971\,
            I => \N__32968\
        );

    \I__6147\ : Span4Mux_v
    port map (
            O => \N__32968\,
            I => \N__32965\
        );

    \I__6146\ : Odrv4
    port map (
            O => \N__32965\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__6145\ : InMux
    port map (
            O => \N__32962\,
            I => \N__32959\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__32959\,
            I => \N__32956\
        );

    \I__6143\ : Odrv12
    port map (
            O => \N__32956\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32950\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__32950\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32944\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__32944\,
            I => \N__32941\
        );

    \I__6138\ : Span4Mux_h
    port map (
            O => \N__32941\,
            I => \N__32938\
        );

    \I__6137\ : Odrv4
    port map (
            O => \N__32938\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32932\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32929\
        );

    \I__6134\ : Span12Mux_h
    port map (
            O => \N__32929\,
            I => \N__32926\
        );

    \I__6133\ : Odrv12
    port map (
            O => \N__32926\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__6132\ : InMux
    port map (
            O => \N__32923\,
            I => \N__32920\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__32920\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32917\,
            I => \N__32914\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__32914\,
            I => \N__32911\
        );

    \I__6128\ : Span4Mux_h
    port map (
            O => \N__32911\,
            I => \N__32908\
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__32908\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32902\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__32902\,
            I => \N__32899\
        );

    \I__6124\ : Span12Mux_s11_v
    port map (
            O => \N__32899\,
            I => \N__32896\
        );

    \I__6123\ : Odrv12
    port map (
            O => \N__32896\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32888\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32885\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32882\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32878\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__32885\,
            I => \N__32873\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__32882\,
            I => \N__32873\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32870\
        );

    \I__6115\ : Span12Mux_v
    port map (
            O => \N__32878\,
            I => \N__32867\
        );

    \I__6114\ : Span12Mux_v
    port map (
            O => \N__32873\,
            I => \N__32864\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32870\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6112\ : Odrv12
    port map (
            O => \N__32867\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6111\ : Odrv12
    port map (
            O => \N__32864\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6110\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32854\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__32854\,
            I => \N__32845\
        );

    \I__6108\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32842\
        );

    \I__6107\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32835\
        );

    \I__6106\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32835\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32835\
        );

    \I__6104\ : CascadeMux
    port map (
            O => \N__32849\,
            I => \N__32832\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32829\
        );

    \I__6102\ : Span4Mux_h
    port map (
            O => \N__32845\,
            I => \N__32814\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__32842\,
            I => \N__32814\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__32835\,
            I => \N__32814\
        );

    \I__6099\ : InMux
    port map (
            O => \N__32832\,
            I => \N__32811\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__32829\,
            I => \N__32808\
        );

    \I__6097\ : InMux
    port map (
            O => \N__32828\,
            I => \N__32805\
        );

    \I__6096\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32790\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32790\
        );

    \I__6094\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32790\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32790\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32790\
        );

    \I__6091\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32790\
        );

    \I__6090\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32790\
        );

    \I__6089\ : Span4Mux_h
    port map (
            O => \N__32814\,
            I => \N__32787\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__32811\,
            I => \N__32778\
        );

    \I__6087\ : Span4Mux_v
    port map (
            O => \N__32808\,
            I => \N__32778\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__32805\,
            I => \N__32778\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__32790\,
            I => \N__32778\
        );

    \I__6084\ : Span4Mux_v
    port map (
            O => \N__32787\,
            I => \N__32775\
        );

    \I__6083\ : Span4Mux_v
    port map (
            O => \N__32778\,
            I => \N__32770\
        );

    \I__6082\ : Span4Mux_v
    port map (
            O => \N__32775\,
            I => \N__32770\
        );

    \I__6081\ : Odrv4
    port map (
            O => \N__32770\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__6080\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32764\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__32764\,
            I => \N__32761\
        );

    \I__6078\ : Span4Mux_h
    port map (
            O => \N__32761\,
            I => \N__32758\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__32758\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32755\,
            I => \N__32752\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__32752\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32746\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__32746\,
            I => \N__32743\
        );

    \I__6072\ : Span4Mux_h
    port map (
            O => \N__32743\,
            I => \N__32740\
        );

    \I__6071\ : Span4Mux_v
    port map (
            O => \N__32740\,
            I => \N__32737\
        );

    \I__6070\ : Odrv4
    port map (
            O => \N__32737\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__6069\ : InMux
    port map (
            O => \N__32734\,
            I => \N__32731\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__32731\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__6067\ : CascadeMux
    port map (
            O => \N__32728\,
            I => \N__32712\
        );

    \I__6066\ : CascadeMux
    port map (
            O => \N__32727\,
            I => \N__32708\
        );

    \I__6065\ : CascadeMux
    port map (
            O => \N__32726\,
            I => \N__32705\
        );

    \I__6064\ : CascadeMux
    port map (
            O => \N__32725\,
            I => \N__32702\
        );

    \I__6063\ : CascadeMux
    port map (
            O => \N__32724\,
            I => \N__32697\
        );

    \I__6062\ : CascadeMux
    port map (
            O => \N__32723\,
            I => \N__32694\
        );

    \I__6061\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32678\
        );

    \I__6060\ : InMux
    port map (
            O => \N__32721\,
            I => \N__32678\
        );

    \I__6059\ : InMux
    port map (
            O => \N__32720\,
            I => \N__32678\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32719\,
            I => \N__32678\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32678\
        );

    \I__6056\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32678\
        );

    \I__6055\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32678\
        );

    \I__6054\ : CascadeMux
    port map (
            O => \N__32715\,
            I => \N__32674\
        );

    \I__6053\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32662\
        );

    \I__6052\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32662\
        );

    \I__6051\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32655\
        );

    \I__6050\ : InMux
    port map (
            O => \N__32705\,
            I => \N__32655\
        );

    \I__6049\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32655\
        );

    \I__6048\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32622\
        );

    \I__6047\ : InMux
    port map (
            O => \N__32700\,
            I => \N__32622\
        );

    \I__6046\ : InMux
    port map (
            O => \N__32697\,
            I => \N__32622\
        );

    \I__6045\ : InMux
    port map (
            O => \N__32694\,
            I => \N__32622\
        );

    \I__6044\ : InMux
    port map (
            O => \N__32693\,
            I => \N__32622\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__32678\,
            I => \N__32619\
        );

    \I__6042\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32610\
        );

    \I__6041\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32610\
        );

    \I__6040\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32610\
        );

    \I__6039\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32610\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__32671\,
            I => \N__32607\
        );

    \I__6037\ : CascadeMux
    port map (
            O => \N__32670\,
            I => \N__32603\
        );

    \I__6036\ : CascadeMux
    port map (
            O => \N__32669\,
            I => \N__32599\
        );

    \I__6035\ : CascadeMux
    port map (
            O => \N__32668\,
            I => \N__32589\
        );

    \I__6034\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32582\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__32662\,
            I => \N__32579\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__32655\,
            I => \N__32576\
        );

    \I__6031\ : CascadeMux
    port map (
            O => \N__32654\,
            I => \N__32573\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__32653\,
            I => \N__32566\
        );

    \I__6029\ : CascadeMux
    port map (
            O => \N__32652\,
            I => \N__32562\
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__32651\,
            I => \N__32558\
        );

    \I__6027\ : CascadeMux
    port map (
            O => \N__32650\,
            I => \N__32554\
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__32649\,
            I => \N__32550\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__32648\,
            I => \N__32546\
        );

    \I__6024\ : CascadeMux
    port map (
            O => \N__32647\,
            I => \N__32542\
        );

    \I__6023\ : CascadeMux
    port map (
            O => \N__32646\,
            I => \N__32538\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32507\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32507\
        );

    \I__6020\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32507\
        );

    \I__6019\ : InMux
    port map (
            O => \N__32642\,
            I => \N__32507\
        );

    \I__6018\ : InMux
    port map (
            O => \N__32641\,
            I => \N__32507\
        );

    \I__6017\ : InMux
    port map (
            O => \N__32640\,
            I => \N__32507\
        );

    \I__6016\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32507\
        );

    \I__6015\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32494\
        );

    \I__6014\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32494\
        );

    \I__6013\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32494\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32494\
        );

    \I__6011\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32494\
        );

    \I__6010\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32494\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__32622\,
            I => \N__32487\
        );

    \I__6008\ : Span4Mux_v
    port map (
            O => \N__32619\,
            I => \N__32487\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__32610\,
            I => \N__32487\
        );

    \I__6006\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32474\
        );

    \I__6005\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32474\
        );

    \I__6004\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32474\
        );

    \I__6003\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32474\
        );

    \I__6002\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32474\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32474\
        );

    \I__6000\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32461\
        );

    \I__5999\ : InMux
    port map (
            O => \N__32596\,
            I => \N__32461\
        );

    \I__5998\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32461\
        );

    \I__5997\ : InMux
    port map (
            O => \N__32594\,
            I => \N__32461\
        );

    \I__5996\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32461\
        );

    \I__5995\ : InMux
    port map (
            O => \N__32592\,
            I => \N__32461\
        );

    \I__5994\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32458\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__32588\,
            I => \N__32448\
        );

    \I__5992\ : CascadeMux
    port map (
            O => \N__32587\,
            I => \N__32440\
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__32586\,
            I => \N__32436\
        );

    \I__5990\ : CascadeMux
    port map (
            O => \N__32585\,
            I => \N__32432\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__32582\,
            I => \N__32428\
        );

    \I__5988\ : Span4Mux_v
    port map (
            O => \N__32579\,
            I => \N__32423\
        );

    \I__5987\ : Span4Mux_v
    port map (
            O => \N__32576\,
            I => \N__32423\
        );

    \I__5986\ : InMux
    port map (
            O => \N__32573\,
            I => \N__32410\
        );

    \I__5985\ : InMux
    port map (
            O => \N__32572\,
            I => \N__32410\
        );

    \I__5984\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32410\
        );

    \I__5983\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32410\
        );

    \I__5982\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32410\
        );

    \I__5981\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32410\
        );

    \I__5980\ : InMux
    port map (
            O => \N__32565\,
            I => \N__32395\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32395\
        );

    \I__5978\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32395\
        );

    \I__5977\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32395\
        );

    \I__5976\ : InMux
    port map (
            O => \N__32557\,
            I => \N__32395\
        );

    \I__5975\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32395\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32553\,
            I => \N__32395\
        );

    \I__5973\ : InMux
    port map (
            O => \N__32550\,
            I => \N__32378\
        );

    \I__5972\ : InMux
    port map (
            O => \N__32549\,
            I => \N__32378\
        );

    \I__5971\ : InMux
    port map (
            O => \N__32546\,
            I => \N__32378\
        );

    \I__5970\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32378\
        );

    \I__5969\ : InMux
    port map (
            O => \N__32542\,
            I => \N__32378\
        );

    \I__5968\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32378\
        );

    \I__5967\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32378\
        );

    \I__5966\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32378\
        );

    \I__5965\ : CascadeMux
    port map (
            O => \N__32536\,
            I => \N__32375\
        );

    \I__5964\ : CascadeMux
    port map (
            O => \N__32535\,
            I => \N__32371\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__32534\,
            I => \N__32367\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__32533\,
            I => \N__32363\
        );

    \I__5961\ : CascadeMux
    port map (
            O => \N__32532\,
            I => \N__32359\
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__32531\,
            I => \N__32355\
        );

    \I__5959\ : CascadeMux
    port map (
            O => \N__32530\,
            I => \N__32351\
        );

    \I__5958\ : CascadeMux
    port map (
            O => \N__32529\,
            I => \N__32347\
        );

    \I__5957\ : CascadeMux
    port map (
            O => \N__32528\,
            I => \N__32343\
        );

    \I__5956\ : CascadeMux
    port map (
            O => \N__32527\,
            I => \N__32339\
        );

    \I__5955\ : CascadeMux
    port map (
            O => \N__32526\,
            I => \N__32335\
        );

    \I__5954\ : CascadeMux
    port map (
            O => \N__32525\,
            I => \N__32331\
        );

    \I__5953\ : CascadeMux
    port map (
            O => \N__32524\,
            I => \N__32327\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__32523\,
            I => \N__32323\
        );

    \I__5951\ : CascadeMux
    port map (
            O => \N__32522\,
            I => \N__32319\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__32507\,
            I => \N__32309\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__32494\,
            I => \N__32309\
        );

    \I__5948\ : Span4Mux_v
    port map (
            O => \N__32487\,
            I => \N__32309\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__32474\,
            I => \N__32309\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__32461\,
            I => \N__32306\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__32458\,
            I => \N__32303\
        );

    \I__5944\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32288\
        );

    \I__5943\ : InMux
    port map (
            O => \N__32456\,
            I => \N__32288\
        );

    \I__5942\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32288\
        );

    \I__5941\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32288\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32288\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32452\,
            I => \N__32288\
        );

    \I__5938\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32288\
        );

    \I__5937\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32281\
        );

    \I__5936\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32281\
        );

    \I__5935\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32281\
        );

    \I__5934\ : InMux
    port map (
            O => \N__32445\,
            I => \N__32278\
        );

    \I__5933\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32261\
        );

    \I__5932\ : InMux
    port map (
            O => \N__32443\,
            I => \N__32261\
        );

    \I__5931\ : InMux
    port map (
            O => \N__32440\,
            I => \N__32261\
        );

    \I__5930\ : InMux
    port map (
            O => \N__32439\,
            I => \N__32261\
        );

    \I__5929\ : InMux
    port map (
            O => \N__32436\,
            I => \N__32261\
        );

    \I__5928\ : InMux
    port map (
            O => \N__32435\,
            I => \N__32261\
        );

    \I__5927\ : InMux
    port map (
            O => \N__32432\,
            I => \N__32261\
        );

    \I__5926\ : InMux
    port map (
            O => \N__32431\,
            I => \N__32261\
        );

    \I__5925\ : Span4Mux_h
    port map (
            O => \N__32428\,
            I => \N__32250\
        );

    \I__5924\ : Span4Mux_h
    port map (
            O => \N__32423\,
            I => \N__32250\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__32410\,
            I => \N__32250\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__32395\,
            I => \N__32250\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32378\,
            I => \N__32250\
        );

    \I__5920\ : InMux
    port map (
            O => \N__32375\,
            I => \N__32233\
        );

    \I__5919\ : InMux
    port map (
            O => \N__32374\,
            I => \N__32233\
        );

    \I__5918\ : InMux
    port map (
            O => \N__32371\,
            I => \N__32233\
        );

    \I__5917\ : InMux
    port map (
            O => \N__32370\,
            I => \N__32233\
        );

    \I__5916\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32233\
        );

    \I__5915\ : InMux
    port map (
            O => \N__32366\,
            I => \N__32233\
        );

    \I__5914\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32233\
        );

    \I__5913\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32233\
        );

    \I__5912\ : InMux
    port map (
            O => \N__32359\,
            I => \N__32216\
        );

    \I__5911\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32216\
        );

    \I__5910\ : InMux
    port map (
            O => \N__32355\,
            I => \N__32216\
        );

    \I__5909\ : InMux
    port map (
            O => \N__32354\,
            I => \N__32216\
        );

    \I__5908\ : InMux
    port map (
            O => \N__32351\,
            I => \N__32216\
        );

    \I__5907\ : InMux
    port map (
            O => \N__32350\,
            I => \N__32216\
        );

    \I__5906\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32216\
        );

    \I__5905\ : InMux
    port map (
            O => \N__32346\,
            I => \N__32216\
        );

    \I__5904\ : InMux
    port map (
            O => \N__32343\,
            I => \N__32199\
        );

    \I__5903\ : InMux
    port map (
            O => \N__32342\,
            I => \N__32199\
        );

    \I__5902\ : InMux
    port map (
            O => \N__32339\,
            I => \N__32199\
        );

    \I__5901\ : InMux
    port map (
            O => \N__32338\,
            I => \N__32199\
        );

    \I__5900\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32199\
        );

    \I__5899\ : InMux
    port map (
            O => \N__32334\,
            I => \N__32199\
        );

    \I__5898\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32199\
        );

    \I__5897\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32199\
        );

    \I__5896\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32186\
        );

    \I__5895\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32186\
        );

    \I__5894\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32186\
        );

    \I__5893\ : InMux
    port map (
            O => \N__32322\,
            I => \N__32186\
        );

    \I__5892\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32186\
        );

    \I__5891\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32186\
        );

    \I__5890\ : Span4Mux_v
    port map (
            O => \N__32309\,
            I => \N__32183\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__32306\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__32303\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__32288\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__32281\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__32278\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__32261\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5883\ : Odrv4
    port map (
            O => \N__32250\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__32233\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__32216\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__32199\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__32186\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5878\ : Odrv4
    port map (
            O => \N__32183\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__5877\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32148\
        );

    \I__5876\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32148\
        );

    \I__5875\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32148\
        );

    \I__5874\ : CascadeMux
    port map (
            O => \N__32155\,
            I => \N__32143\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__32148\,
            I => \N__32129\
        );

    \I__5872\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32125\
        );

    \I__5871\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32096\
        );

    \I__5870\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32096\
        );

    \I__5869\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32096\
        );

    \I__5868\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32096\
        );

    \I__5867\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32096\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__32139\,
            I => \N__32093\
        );

    \I__5865\ : InMux
    port map (
            O => \N__32138\,
            I => \N__32083\
        );

    \I__5864\ : InMux
    port map (
            O => \N__32137\,
            I => \N__32070\
        );

    \I__5863\ : InMux
    port map (
            O => \N__32136\,
            I => \N__32070\
        );

    \I__5862\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32070\
        );

    \I__5861\ : InMux
    port map (
            O => \N__32134\,
            I => \N__32070\
        );

    \I__5860\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32070\
        );

    \I__5859\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32070\
        );

    \I__5858\ : Span4Mux_v
    port map (
            O => \N__32129\,
            I => \N__32067\
        );

    \I__5857\ : InMux
    port map (
            O => \N__32128\,
            I => \N__32064\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__32125\,
            I => \N__32061\
        );

    \I__5855\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32050\
        );

    \I__5854\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32050\
        );

    \I__5853\ : InMux
    port map (
            O => \N__32122\,
            I => \N__32050\
        );

    \I__5852\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32050\
        );

    \I__5851\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32050\
        );

    \I__5850\ : InMux
    port map (
            O => \N__32119\,
            I => \N__32037\
        );

    \I__5849\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32037\
        );

    \I__5848\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32037\
        );

    \I__5847\ : InMux
    port map (
            O => \N__32116\,
            I => \N__32037\
        );

    \I__5846\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32037\
        );

    \I__5845\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32037\
        );

    \I__5844\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32026\
        );

    \I__5843\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32026\
        );

    \I__5842\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32026\
        );

    \I__5841\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32026\
        );

    \I__5840\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32026\
        );

    \I__5839\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32022\
        );

    \I__5838\ : CascadeMux
    port map (
            O => \N__32107\,
            I => \N__32019\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__32096\,
            I => \N__32011\
        );

    \I__5836\ : InMux
    port map (
            O => \N__32093\,
            I => \N__31994\
        );

    \I__5835\ : InMux
    port map (
            O => \N__32092\,
            I => \N__31994\
        );

    \I__5834\ : InMux
    port map (
            O => \N__32091\,
            I => \N__31994\
        );

    \I__5833\ : InMux
    port map (
            O => \N__32090\,
            I => \N__31994\
        );

    \I__5832\ : InMux
    port map (
            O => \N__32089\,
            I => \N__31994\
        );

    \I__5831\ : InMux
    port map (
            O => \N__32088\,
            I => \N__31994\
        );

    \I__5830\ : InMux
    port map (
            O => \N__32087\,
            I => \N__31994\
        );

    \I__5829\ : InMux
    port map (
            O => \N__32086\,
            I => \N__31994\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__32083\,
            I => \N__31982\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__32070\,
            I => \N__31977\
        );

    \I__5826\ : Span4Mux_h
    port map (
            O => \N__32067\,
            I => \N__31977\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__32064\,
            I => \N__31968\
        );

    \I__5824\ : Span4Mux_v
    port map (
            O => \N__32061\,
            I => \N__31968\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__32050\,
            I => \N__31968\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__31968\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__32026\,
            I => \N__31965\
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__32025\,
            I => \N__31953\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__32022\,
            I => \N__31946\
        );

    \I__5818\ : InMux
    port map (
            O => \N__32019\,
            I => \N__31933\
        );

    \I__5817\ : InMux
    port map (
            O => \N__32018\,
            I => \N__31933\
        );

    \I__5816\ : InMux
    port map (
            O => \N__32017\,
            I => \N__31933\
        );

    \I__5815\ : InMux
    port map (
            O => \N__32016\,
            I => \N__31933\
        );

    \I__5814\ : InMux
    port map (
            O => \N__32015\,
            I => \N__31933\
        );

    \I__5813\ : InMux
    port map (
            O => \N__32014\,
            I => \N__31933\
        );

    \I__5812\ : Span4Mux_v
    port map (
            O => \N__32011\,
            I => \N__31928\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__31994\,
            I => \N__31928\
        );

    \I__5810\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31913\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31913\
        );

    \I__5808\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31913\
        );

    \I__5807\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31913\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31913\
        );

    \I__5805\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31913\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31913\
        );

    \I__5803\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31908\
        );

    \I__5802\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31908\
        );

    \I__5801\ : Span12Mux_s11_h
    port map (
            O => \N__31982\,
            I => \N__31905\
        );

    \I__5800\ : Span4Mux_v
    port map (
            O => \N__31977\,
            I => \N__31902\
        );

    \I__5799\ : Span4Mux_v
    port map (
            O => \N__31968\,
            I => \N__31897\
        );

    \I__5798\ : Span4Mux_v
    port map (
            O => \N__31965\,
            I => \N__31897\
        );

    \I__5797\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31882\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31882\
        );

    \I__5795\ : InMux
    port map (
            O => \N__31962\,
            I => \N__31882\
        );

    \I__5794\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31882\
        );

    \I__5793\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31882\
        );

    \I__5792\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31882\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31882\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31879\
        );

    \I__5789\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31866\
        );

    \I__5788\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31866\
        );

    \I__5787\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31866\
        );

    \I__5786\ : InMux
    port map (
            O => \N__31951\,
            I => \N__31866\
        );

    \I__5785\ : InMux
    port map (
            O => \N__31950\,
            I => \N__31866\
        );

    \I__5784\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31866\
        );

    \I__5783\ : Span4Mux_h
    port map (
            O => \N__31946\,
            I => \N__31859\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__31933\,
            I => \N__31859\
        );

    \I__5781\ : Span4Mux_h
    port map (
            O => \N__31928\,
            I => \N__31859\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31913\,
            I => \N__31854\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__31908\,
            I => \N__31854\
        );

    \I__5778\ : Odrv12
    port map (
            O => \N__31905\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5777\ : Odrv4
    port map (
            O => \N__31902\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__31897\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__31882\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__31879\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__31866\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__31859\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5771\ : Odrv12
    port map (
            O => \N__31854\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5770\ : CascadeMux
    port map (
            O => \N__31837\,
            I => \N__31834\
        );

    \I__5769\ : InMux
    port map (
            O => \N__31834\,
            I => \N__31831\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__31831\,
            I => \N__31826\
        );

    \I__5767\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31823\
        );

    \I__5766\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31820\
        );

    \I__5765\ : Span12Mux_h
    port map (
            O => \N__31826\,
            I => \N__31817\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__31823\,
            I => \N__31814\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__31820\,
            I => \N__31811\
        );

    \I__5762\ : Odrv12
    port map (
            O => \N__31817\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__5761\ : Odrv12
    port map (
            O => \N__31814\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__31811\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__31804\,
            I => \N__31800\
        );

    \I__5758\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31797\
        );

    \I__5757\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31794\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__31797\,
            I => \N__31789\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__31794\,
            I => \N__31789\
        );

    \I__5754\ : Span4Mux_v
    port map (
            O => \N__31789\,
            I => \N__31785\
        );

    \I__5753\ : CascadeMux
    port map (
            O => \N__31788\,
            I => \N__31782\
        );

    \I__5752\ : Span4Mux_h
    port map (
            O => \N__31785\,
            I => \N__31778\
        );

    \I__5751\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31775\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31772\
        );

    \I__5749\ : Span4Mux_h
    port map (
            O => \N__31778\,
            I => \N__31767\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__31775\,
            I => \N__31767\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__31772\,
            I => \N__31764\
        );

    \I__5746\ : Odrv4
    port map (
            O => \N__31767\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__5745\ : Odrv4
    port map (
            O => \N__31764\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__5744\ : InMux
    port map (
            O => \N__31759\,
            I => \N__31756\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__31756\,
            I => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__31753\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_\
        );

    \I__5741\ : CascadeMux
    port map (
            O => \N__31750\,
            I => \elapsed_time_ns_1_RNIRB3CP1_0_3_cascade_\
        );

    \I__5740\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31744\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__31744\,
            I => \N__31741\
        );

    \I__5738\ : Span4Mux_v
    port map (
            O => \N__31741\,
            I => \N__31738\
        );

    \I__5737\ : Odrv4
    port map (
            O => \N__31738\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__5736\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31732\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__31732\,
            I => \N__31729\
        );

    \I__5734\ : Odrv4
    port map (
            O => \N__31729\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__5733\ : CascadeMux
    port map (
            O => \N__31726\,
            I => \N__31723\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31720\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__31720\,
            I => \N__31717\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__31717\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__31714\,
            I => \N__31711\
        );

    \I__5728\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31708\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__31708\,
            I => \N__31705\
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__31705\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__5725\ : InMux
    port map (
            O => \N__31702\,
            I => \N__31699\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__31699\,
            I => \N__31696\
        );

    \I__5723\ : Odrv4
    port map (
            O => \N__31696\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__5722\ : InMux
    port map (
            O => \N__31693\,
            I => \N__31690\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__31690\,
            I => \N__31687\
        );

    \I__5720\ : Span4Mux_v
    port map (
            O => \N__31687\,
            I => \N__31684\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__31684\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__5718\ : InMux
    port map (
            O => \N__31681\,
            I => \N__31678\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__31678\,
            I => \N__31675\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__31675\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__5715\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31669\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__31669\,
            I => \N__31666\
        );

    \I__5713\ : Span4Mux_h
    port map (
            O => \N__31666\,
            I => \N__31663\
        );

    \I__5712\ : Span4Mux_v
    port map (
            O => \N__31663\,
            I => \N__31660\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__31660\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__5710\ : InMux
    port map (
            O => \N__31657\,
            I => \N__31654\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__31654\,
            I => \N__31649\
        );

    \I__5708\ : InMux
    port map (
            O => \N__31653\,
            I => \N__31646\
        );

    \I__5707\ : InMux
    port map (
            O => \N__31652\,
            I => \N__31643\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__31649\,
            I => \N__31639\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__31646\,
            I => \N__31636\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__31643\,
            I => \N__31633\
        );

    \I__5703\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31630\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__31639\,
            I => \N__31627\
        );

    \I__5701\ : Span4Mux_h
    port map (
            O => \N__31636\,
            I => \N__31624\
        );

    \I__5700\ : Span12Mux_h
    port map (
            O => \N__31633\,
            I => \N__31619\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__31630\,
            I => \N__31619\
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__31627\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__31624\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5696\ : Odrv12
    port map (
            O => \N__31619\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__5695\ : CascadeMux
    port map (
            O => \N__31612\,
            I => \N__31609\
        );

    \I__5694\ : InMux
    port map (
            O => \N__31609\,
            I => \N__31605\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__31608\,
            I => \N__31602\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__31605\,
            I => \N__31599\
        );

    \I__5691\ : InMux
    port map (
            O => \N__31602\,
            I => \N__31596\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__31599\,
            I => \N__31590\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__31596\,
            I => \N__31590\
        );

    \I__5688\ : InMux
    port map (
            O => \N__31595\,
            I => \N__31587\
        );

    \I__5687\ : Span4Mux_h
    port map (
            O => \N__31590\,
            I => \N__31584\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__31587\,
            I => \N__31581\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__31584\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__5684\ : Odrv12
    port map (
            O => \N__31581\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__31576\,
            I => \N__31573\
        );

    \I__5682\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31570\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__31570\,
            I => \N__31567\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__31567\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__5679\ : CascadeMux
    port map (
            O => \N__31564\,
            I => \N__31560\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__31563\,
            I => \N__31557\
        );

    \I__5677\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31554\
        );

    \I__5676\ : InMux
    port map (
            O => \N__31557\,
            I => \N__31551\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__31554\,
            I => \N__31548\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__31551\,
            I => \N__31545\
        );

    \I__5673\ : Span4Mux_h
    port map (
            O => \N__31548\,
            I => \N__31540\
        );

    \I__5672\ : Span4Mux_h
    port map (
            O => \N__31545\,
            I => \N__31537\
        );

    \I__5671\ : InMux
    port map (
            O => \N__31544\,
            I => \N__31534\
        );

    \I__5670\ : InMux
    port map (
            O => \N__31543\,
            I => \N__31531\
        );

    \I__5669\ : Span4Mux_v
    port map (
            O => \N__31540\,
            I => \N__31528\
        );

    \I__5668\ : Span4Mux_h
    port map (
            O => \N__31537\,
            I => \N__31521\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__31534\,
            I => \N__31521\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__31531\,
            I => \N__31521\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__31528\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__5664\ : Odrv4
    port map (
            O => \N__31521\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__5663\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31513\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__31513\,
            I => \N__31509\
        );

    \I__5661\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31505\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__31509\,
            I => \N__31502\
        );

    \I__5659\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31499\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__31505\,
            I => \N__31496\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__31502\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__31499\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__5655\ : Odrv12
    port map (
            O => \N__31496\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__5654\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31486\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__31486\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__5652\ : InMux
    port map (
            O => \N__31483\,
            I => \N__31480\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__31480\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__5650\ : InMux
    port map (
            O => \N__31477\,
            I => \N__31474\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__31474\,
            I => \N__31471\
        );

    \I__5648\ : Span4Mux_v
    port map (
            O => \N__31471\,
            I => \N__31468\
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__31468\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__5646\ : InMux
    port map (
            O => \N__31465\,
            I => \N__31462\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__31462\,
            I => \N__31459\
        );

    \I__5644\ : Odrv12
    port map (
            O => \N__31459\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__31456\,
            I => \N__31453\
        );

    \I__5642\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31450\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__31450\,
            I => \N__31446\
        );

    \I__5640\ : InMux
    port map (
            O => \N__31449\,
            I => \N__31443\
        );

    \I__5639\ : Span4Mux_v
    port map (
            O => \N__31446\,
            I => \N__31439\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__31443\,
            I => \N__31436\
        );

    \I__5637\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31433\
        );

    \I__5636\ : Span4Mux_h
    port map (
            O => \N__31439\,
            I => \N__31428\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__31436\,
            I => \N__31428\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__31433\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5633\ : Odrv4
    port map (
            O => \N__31428\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5632\ : CascadeMux
    port map (
            O => \N__31423\,
            I => \N__31420\
        );

    \I__5631\ : InMux
    port map (
            O => \N__31420\,
            I => \N__31416\
        );

    \I__5630\ : InMux
    port map (
            O => \N__31419\,
            I => \N__31413\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__31416\,
            I => \N__31410\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__31413\,
            I => \N__31407\
        );

    \I__5627\ : Span4Mux_h
    port map (
            O => \N__31410\,
            I => \N__31403\
        );

    \I__5626\ : Span4Mux_v
    port map (
            O => \N__31407\,
            I => \N__31400\
        );

    \I__5625\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31397\
        );

    \I__5624\ : Span4Mux_v
    port map (
            O => \N__31403\,
            I => \N__31393\
        );

    \I__5623\ : Span4Mux_h
    port map (
            O => \N__31400\,
            I => \N__31388\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31388\
        );

    \I__5621\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31385\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__31393\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__31388\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__31385\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__31378\,
            I => \N__31375\
        );

    \I__5616\ : InMux
    port map (
            O => \N__31375\,
            I => \N__31372\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__31372\,
            I => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__31369\,
            I => \N__31365\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__31368\,
            I => \N__31362\
        );

    \I__5612\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31359\
        );

    \I__5611\ : InMux
    port map (
            O => \N__31362\,
            I => \N__31356\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__31359\,
            I => \N__31353\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__31356\,
            I => \N__31348\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__31353\,
            I => \N__31345\
        );

    \I__5607\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31342\
        );

    \I__5606\ : InMux
    port map (
            O => \N__31351\,
            I => \N__31339\
        );

    \I__5605\ : Span4Mux_v
    port map (
            O => \N__31348\,
            I => \N__31336\
        );

    \I__5604\ : Span4Mux_v
    port map (
            O => \N__31345\,
            I => \N__31331\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__31342\,
            I => \N__31331\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__31339\,
            I => \N__31328\
        );

    \I__5601\ : Span4Mux_h
    port map (
            O => \N__31336\,
            I => \N__31325\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__31331\,
            I => \N__31322\
        );

    \I__5599\ : Span4Mux_v
    port map (
            O => \N__31328\,
            I => \N__31319\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__31325\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__31322\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__5596\ : Odrv4
    port map (
            O => \N__31319\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__5595\ : InMux
    port map (
            O => \N__31312\,
            I => \N__31308\
        );

    \I__5594\ : InMux
    port map (
            O => \N__31311\,
            I => \N__31305\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__31308\,
            I => \N__31302\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__31305\,
            I => \N__31298\
        );

    \I__5591\ : Span4Mux_h
    port map (
            O => \N__31302\,
            I => \N__31295\
        );

    \I__5590\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31292\
        );

    \I__5589\ : Span4Mux_v
    port map (
            O => \N__31298\,
            I => \N__31289\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__31295\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__31292\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__31289\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__5585\ : CascadeMux
    port map (
            O => \N__31282\,
            I => \N__31279\
        );

    \I__5584\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31276\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__31276\,
            I => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\
        );

    \I__5582\ : CascadeMux
    port map (
            O => \N__31273\,
            I => \N__31270\
        );

    \I__5581\ : InMux
    port map (
            O => \N__31270\,
            I => \N__31267\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__31267\,
            I => \N__31263\
        );

    \I__5579\ : InMux
    port map (
            O => \N__31266\,
            I => \N__31259\
        );

    \I__5578\ : Span4Mux_h
    port map (
            O => \N__31263\,
            I => \N__31256\
        );

    \I__5577\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31253\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__31259\,
            I => \N__31250\
        );

    \I__5575\ : Odrv4
    port map (
            O => \N__31256\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__31253\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__31250\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__31243\,
            I => \N__31240\
        );

    \I__5571\ : InMux
    port map (
            O => \N__31240\,
            I => \N__31236\
        );

    \I__5570\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31233\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__31236\,
            I => \N__31229\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__31233\,
            I => \N__31225\
        );

    \I__5567\ : InMux
    port map (
            O => \N__31232\,
            I => \N__31222\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__31229\,
            I => \N__31219\
        );

    \I__5565\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31216\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__31225\,
            I => \N__31211\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__31222\,
            I => \N__31211\
        );

    \I__5562\ : Span4Mux_v
    port map (
            O => \N__31219\,
            I => \N__31208\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__31216\,
            I => \N__31203\
        );

    \I__5560\ : Span4Mux_h
    port map (
            O => \N__31211\,
            I => \N__31203\
        );

    \I__5559\ : Odrv4
    port map (
            O => \N__31208\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__5558\ : Odrv4
    port map (
            O => \N__31203\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__5557\ : CascadeMux
    port map (
            O => \N__31198\,
            I => \N__31195\
        );

    \I__5556\ : InMux
    port map (
            O => \N__31195\,
            I => \N__31192\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__31192\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__5554\ : CascadeMux
    port map (
            O => \N__31189\,
            I => \N__31186\
        );

    \I__5553\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31183\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31179\
        );

    \I__5551\ : InMux
    port map (
            O => \N__31182\,
            I => \N__31176\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__31179\,
            I => \N__31173\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__31176\,
            I => \N__31170\
        );

    \I__5548\ : Span4Mux_v
    port map (
            O => \N__31173\,
            I => \N__31165\
        );

    \I__5547\ : Span4Mux_h
    port map (
            O => \N__31170\,
            I => \N__31162\
        );

    \I__5546\ : InMux
    port map (
            O => \N__31169\,
            I => \N__31159\
        );

    \I__5545\ : InMux
    port map (
            O => \N__31168\,
            I => \N__31156\
        );

    \I__5544\ : Span4Mux_h
    port map (
            O => \N__31165\,
            I => \N__31153\
        );

    \I__5543\ : Span4Mux_h
    port map (
            O => \N__31162\,
            I => \N__31150\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__31159\,
            I => \N__31145\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__31156\,
            I => \N__31145\
        );

    \I__5540\ : Odrv4
    port map (
            O => \N__31153\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__5539\ : Odrv4
    port map (
            O => \N__31150\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__5538\ : Odrv12
    port map (
            O => \N__31145\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__5537\ : InMux
    port map (
            O => \N__31138\,
            I => \N__31134\
        );

    \I__5536\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31131\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31127\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__31131\,
            I => \N__31124\
        );

    \I__5533\ : InMux
    port map (
            O => \N__31130\,
            I => \N__31121\
        );

    \I__5532\ : Span4Mux_h
    port map (
            O => \N__31127\,
            I => \N__31116\
        );

    \I__5531\ : Span4Mux_v
    port map (
            O => \N__31124\,
            I => \N__31116\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__31121\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__5529\ : Odrv4
    port map (
            O => \N__31116\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__5528\ : CascadeMux
    port map (
            O => \N__31111\,
            I => \N__31108\
        );

    \I__5527\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31105\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__31105\,
            I => \N__31102\
        );

    \I__5525\ : Odrv12
    port map (
            O => \N__31102\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__5524\ : CascadeMux
    port map (
            O => \N__31099\,
            I => \N__31096\
        );

    \I__5523\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31092\
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__31095\,
            I => \N__31089\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__31092\,
            I => \N__31085\
        );

    \I__5520\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31082\
        );

    \I__5519\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31079\
        );

    \I__5518\ : Span4Mux_h
    port map (
            O => \N__31085\,
            I => \N__31076\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__31082\,
            I => \N__31073\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__31079\,
            I => \N__31070\
        );

    \I__5515\ : Odrv4
    port map (
            O => \N__31076\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__5514\ : Odrv12
    port map (
            O => \N__31073\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__5513\ : Odrv12
    port map (
            O => \N__31070\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__5512\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31060\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__31060\,
            I => \N__31055\
        );

    \I__5510\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31052\
        );

    \I__5509\ : InMux
    port map (
            O => \N__31058\,
            I => \N__31049\
        );

    \I__5508\ : Span4Mux_v
    port map (
            O => \N__31055\,
            I => \N__31043\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__31052\,
            I => \N__31043\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__31049\,
            I => \N__31040\
        );

    \I__5505\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31037\
        );

    \I__5504\ : Span4Mux_h
    port map (
            O => \N__31043\,
            I => \N__31034\
        );

    \I__5503\ : Span12Mux_h
    port map (
            O => \N__31040\,
            I => \N__31029\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__31037\,
            I => \N__31029\
        );

    \I__5501\ : Odrv4
    port map (
            O => \N__31034\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__5500\ : Odrv12
    port map (
            O => \N__31029\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__5499\ : InMux
    port map (
            O => \N__31024\,
            I => \N__31021\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__31021\,
            I => \N__31018\
        );

    \I__5497\ : Odrv12
    port map (
            O => \N__31018\,
            I => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\
        );

    \I__5496\ : CascadeMux
    port map (
            O => \N__31015\,
            I => \N__31011\
        );

    \I__5495\ : CascadeMux
    port map (
            O => \N__31014\,
            I => \N__31008\
        );

    \I__5494\ : InMux
    port map (
            O => \N__31011\,
            I => \N__31005\
        );

    \I__5493\ : InMux
    port map (
            O => \N__31008\,
            I => \N__31002\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__31005\,
            I => \N__30998\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__31002\,
            I => \N__30995\
        );

    \I__5490\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30992\
        );

    \I__5489\ : Span4Mux_h
    port map (
            O => \N__30998\,
            I => \N__30985\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__30995\,
            I => \N__30985\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__30992\,
            I => \N__30985\
        );

    \I__5486\ : Span4Mux_h
    port map (
            O => \N__30985\,
            I => \N__30982\
        );

    \I__5485\ : Span4Mux_v
    port map (
            O => \N__30982\,
            I => \N__30978\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30975\
        );

    \I__5483\ : Odrv4
    port map (
            O => \N__30978\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__30975\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30967\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30967\,
            I => \N__30964\
        );

    \I__5479\ : Span4Mux_h
    port map (
            O => \N__30964\,
            I => \N__30959\
        );

    \I__5478\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30956\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30953\
        );

    \I__5476\ : Odrv4
    port map (
            O => \N__30959\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30956\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__30953\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30943\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__30943\,
            I => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__30940\,
            I => \N__30936\
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__30939\,
            I => \N__30933\
        );

    \I__5469\ : InMux
    port map (
            O => \N__30936\,
            I => \N__30930\
        );

    \I__5468\ : InMux
    port map (
            O => \N__30933\,
            I => \N__30927\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__30930\,
            I => \N__30924\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__30927\,
            I => \N__30920\
        );

    \I__5465\ : Span4Mux_v
    port map (
            O => \N__30924\,
            I => \N__30916\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30923\,
            I => \N__30913\
        );

    \I__5463\ : Span4Mux_h
    port map (
            O => \N__30920\,
            I => \N__30910\
        );

    \I__5462\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30907\
        );

    \I__5461\ : Span4Mux_h
    port map (
            O => \N__30916\,
            I => \N__30902\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__30913\,
            I => \N__30902\
        );

    \I__5459\ : Sp12to4
    port map (
            O => \N__30910\,
            I => \N__30897\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__30907\,
            I => \N__30897\
        );

    \I__5457\ : Odrv4
    port map (
            O => \N__30902\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__5456\ : Odrv12
    port map (
            O => \N__30897\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30889\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__30889\,
            I => \N__30885\
        );

    \I__5453\ : InMux
    port map (
            O => \N__30888\,
            I => \N__30881\
        );

    \I__5452\ : Span4Mux_v
    port map (
            O => \N__30885\,
            I => \N__30878\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30884\,
            I => \N__30875\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__30881\,
            I => \N__30872\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__30878\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__30875\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__5447\ : Odrv12
    port map (
            O => \N__30872\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30865\,
            I => \N__30862\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__30862\,
            I => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\
        );

    \I__5444\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30856\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__30856\,
            I => \N__30853\
        );

    \I__5442\ : Odrv4
    port map (
            O => \N__30853\,
            I => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\
        );

    \I__5441\ : CascadeMux
    port map (
            O => \N__30850\,
            I => \N__30846\
        );

    \I__5440\ : CascadeMux
    port map (
            O => \N__30849\,
            I => \N__30843\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30840\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30837\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__30840\,
            I => \N__30834\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__30837\,
            I => \N__30831\
        );

    \I__5435\ : Span4Mux_h
    port map (
            O => \N__30834\,
            I => \N__30826\
        );

    \I__5434\ : Span4Mux_v
    port map (
            O => \N__30831\,
            I => \N__30823\
        );

    \I__5433\ : InMux
    port map (
            O => \N__30830\,
            I => \N__30820\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30817\
        );

    \I__5431\ : Span4Mux_v
    port map (
            O => \N__30826\,
            I => \N__30814\
        );

    \I__5430\ : Span4Mux_h
    port map (
            O => \N__30823\,
            I => \N__30809\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__30820\,
            I => \N__30809\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__30817\,
            I => \N__30806\
        );

    \I__5427\ : Odrv4
    port map (
            O => \N__30814\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__5426\ : Odrv4
    port map (
            O => \N__30809\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__5425\ : Odrv12
    port map (
            O => \N__30806\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__5424\ : InMux
    port map (
            O => \N__30799\,
            I => \N__30795\
        );

    \I__5423\ : InMux
    port map (
            O => \N__30798\,
            I => \N__30792\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__30795\,
            I => \N__30788\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__30792\,
            I => \N__30785\
        );

    \I__5420\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30782\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__30788\,
            I => \N__30777\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__30785\,
            I => \N__30777\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__30782\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__5416\ : Odrv4
    port map (
            O => \N__30777\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__5415\ : InMux
    port map (
            O => \N__30772\,
            I => \N__30769\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__30769\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__5413\ : CascadeMux
    port map (
            O => \N__30766\,
            I => \N__30762\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__30765\,
            I => \N__30759\
        );

    \I__5411\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30756\
        );

    \I__5410\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30753\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30750\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__30753\,
            I => \N__30746\
        );

    \I__5407\ : Span4Mux_h
    port map (
            O => \N__30750\,
            I => \N__30742\
        );

    \I__5406\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30739\
        );

    \I__5405\ : Span4Mux_h
    port map (
            O => \N__30746\,
            I => \N__30736\
        );

    \I__5404\ : InMux
    port map (
            O => \N__30745\,
            I => \N__30733\
        );

    \I__5403\ : Span4Mux_h
    port map (
            O => \N__30742\,
            I => \N__30728\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__30739\,
            I => \N__30728\
        );

    \I__5401\ : Sp12to4
    port map (
            O => \N__30736\,
            I => \N__30723\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__30733\,
            I => \N__30723\
        );

    \I__5399\ : Odrv4
    port map (
            O => \N__30728\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__5398\ : Odrv12
    port map (
            O => \N__30723\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__5397\ : InMux
    port map (
            O => \N__30718\,
            I => \N__30715\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__30715\,
            I => \N__30710\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30714\,
            I => \N__30707\
        );

    \I__5394\ : InMux
    port map (
            O => \N__30713\,
            I => \N__30704\
        );

    \I__5393\ : Span12Mux_v
    port map (
            O => \N__30710\,
            I => \N__30701\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__30707\,
            I => \N__30698\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__30704\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__5390\ : Odrv12
    port map (
            O => \N__30701\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__5389\ : Odrv4
    port map (
            O => \N__30698\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__5388\ : InMux
    port map (
            O => \N__30691\,
            I => \N__30688\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__30688\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__5386\ : CascadeMux
    port map (
            O => \N__30685\,
            I => \N__30682\
        );

    \I__5385\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30676\
        );

    \I__5384\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30676\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__30676\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__5382\ : CascadeMux
    port map (
            O => \N__30673\,
            I => \N__30670\
        );

    \I__5381\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30661\
        );

    \I__5380\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30661\
        );

    \I__5379\ : InMux
    port map (
            O => \N__30668\,
            I => \N__30661\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__30661\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__5377\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30649\
        );

    \I__5376\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30639\
        );

    \I__5375\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30636\
        );

    \I__5374\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30631\
        );

    \I__5373\ : InMux
    port map (
            O => \N__30654\,
            I => \N__30631\
        );

    \I__5372\ : InMux
    port map (
            O => \N__30653\,
            I => \N__30625\
        );

    \I__5371\ : InMux
    port map (
            O => \N__30652\,
            I => \N__30625\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30612\
        );

    \I__5369\ : InMux
    port map (
            O => \N__30648\,
            I => \N__30597\
        );

    \I__5368\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30597\
        );

    \I__5367\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30597\
        );

    \I__5366\ : InMux
    port map (
            O => \N__30645\,
            I => \N__30597\
        );

    \I__5365\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30597\
        );

    \I__5364\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30597\
        );

    \I__5363\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30597\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30592\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__30636\,
            I => \N__30592\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__30631\,
            I => \N__30589\
        );

    \I__5359\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30586\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__30625\,
            I => \N__30583\
        );

    \I__5357\ : InMux
    port map (
            O => \N__30624\,
            I => \N__30578\
        );

    \I__5356\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30578\
        );

    \I__5355\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30573\
        );

    \I__5354\ : InMux
    port map (
            O => \N__30621\,
            I => \N__30573\
        );

    \I__5353\ : InMux
    port map (
            O => \N__30620\,
            I => \N__30570\
        );

    \I__5352\ : InMux
    port map (
            O => \N__30619\,
            I => \N__30559\
        );

    \I__5351\ : InMux
    port map (
            O => \N__30618\,
            I => \N__30559\
        );

    \I__5350\ : InMux
    port map (
            O => \N__30617\,
            I => \N__30559\
        );

    \I__5349\ : InMux
    port map (
            O => \N__30616\,
            I => \N__30559\
        );

    \I__5348\ : InMux
    port map (
            O => \N__30615\,
            I => \N__30559\
        );

    \I__5347\ : Span4Mux_h
    port map (
            O => \N__30612\,
            I => \N__30552\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__30597\,
            I => \N__30552\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__30592\,
            I => \N__30552\
        );

    \I__5344\ : Odrv4
    port map (
            O => \N__30589\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__30586\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__30583\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__30578\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__30573\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__30570\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__30559\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__30552\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__30535\,
            I => \N__30532\
        );

    \I__5335\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30528\
        );

    \I__5334\ : InMux
    port map (
            O => \N__30531\,
            I => \N__30525\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__30528\,
            I => \N__30522\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__30525\,
            I => \N__30519\
        );

    \I__5331\ : Span4Mux_h
    port map (
            O => \N__30522\,
            I => \N__30514\
        );

    \I__5330\ : Span4Mux_h
    port map (
            O => \N__30519\,
            I => \N__30514\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__30514\,
            I => \N__30509\
        );

    \I__5328\ : InMux
    port map (
            O => \N__30513\,
            I => \N__30506\
        );

    \I__5327\ : InMux
    port map (
            O => \N__30512\,
            I => \N__30503\
        );

    \I__5326\ : Span4Mux_h
    port map (
            O => \N__30509\,
            I => \N__30500\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__30506\,
            I => \N__30495\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__30503\,
            I => \N__30495\
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__30500\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__5322\ : Odrv12
    port map (
            O => \N__30495\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__5321\ : InMux
    port map (
            O => \N__30490\,
            I => \N__30487\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__30487\,
            I => \N__30482\
        );

    \I__5319\ : InMux
    port map (
            O => \N__30486\,
            I => \N__30479\
        );

    \I__5318\ : InMux
    port map (
            O => \N__30485\,
            I => \N__30476\
        );

    \I__5317\ : Span4Mux_v
    port map (
            O => \N__30482\,
            I => \N__30473\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__30479\,
            I => \N__30470\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__30476\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__5314\ : Odrv4
    port map (
            O => \N__30473\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__5313\ : Odrv12
    port map (
            O => \N__30470\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__5312\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30460\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__30460\,
            I => \N__30457\
        );

    \I__5310\ : Span4Mux_v
    port map (
            O => \N__30457\,
            I => \N__30454\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__30454\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30448\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__30448\,
            I => \N__30445\
        );

    \I__5306\ : Odrv4
    port map (
            O => \N__30445\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__5305\ : InMux
    port map (
            O => \N__30442\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__5304\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30436\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__30436\,
            I => \N__30433\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__30433\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__5301\ : InMux
    port map (
            O => \N__30430\,
            I => \bfn_12_12_0_\
        );

    \I__5300\ : InMux
    port map (
            O => \N__30427\,
            I => \N__30424\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30421\
        );

    \I__5298\ : Odrv4
    port map (
            O => \N__30421\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__5297\ : InMux
    port map (
            O => \N__30418\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__5296\ : InMux
    port map (
            O => \N__30415\,
            I => \N__30412\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__30412\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__5294\ : InMux
    port map (
            O => \N__30409\,
            I => \N__30406\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__30406\,
            I => \N__30403\
        );

    \I__5292\ : Odrv4
    port map (
            O => \N__30403\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__5291\ : InMux
    port map (
            O => \N__30400\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__5290\ : InMux
    port map (
            O => \N__30397\,
            I => \N__30394\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__30394\,
            I => \N__30391\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__30391\,
            I => \N__30388\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__30388\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__5286\ : InMux
    port map (
            O => \N__30385\,
            I => \N__30382\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__30382\,
            I => \N__30379\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__30379\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30376\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30373\,
            I => \N__30370\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__30370\,
            I => \N__30367\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__30367\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__5279\ : InMux
    port map (
            O => \N__30364\,
            I => \N__30361\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__30361\,
            I => \N__30358\
        );

    \I__5277\ : Odrv4
    port map (
            O => \N__30358\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__5276\ : InMux
    port map (
            O => \N__30355\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__5275\ : InMux
    port map (
            O => \N__30352\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__5274\ : InMux
    port map (
            O => \N__30349\,
            I => \N__30346\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__30346\,
            I => \N__30343\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__30343\,
            I => \current_shift_inst.control_input_31\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__30340\,
            I => \current_shift_inst.control_input_31_cascade_\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30334\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__30334\,
            I => \N__30331\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__30331\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__5267\ : InMux
    port map (
            O => \N__30328\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__5266\ : CascadeMux
    port map (
            O => \N__30325\,
            I => \N__30322\
        );

    \I__5265\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30319\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__30319\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__30316\,
            I => \N__30313\
        );

    \I__5262\ : InMux
    port map (
            O => \N__30313\,
            I => \N__30308\
        );

    \I__5261\ : InMux
    port map (
            O => \N__30312\,
            I => \N__30305\
        );

    \I__5260\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30301\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__30308\,
            I => \N__30298\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__30305\,
            I => \N__30295\
        );

    \I__5257\ : InMux
    port map (
            O => \N__30304\,
            I => \N__30292\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__30301\,
            I => \N__30288\
        );

    \I__5255\ : Span4Mux_v
    port map (
            O => \N__30298\,
            I => \N__30281\
        );

    \I__5254\ : Span4Mux_h
    port map (
            O => \N__30295\,
            I => \N__30281\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__30292\,
            I => \N__30281\
        );

    \I__5252\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30278\
        );

    \I__5251\ : Span4Mux_v
    port map (
            O => \N__30288\,
            I => \N__30273\
        );

    \I__5250\ : Span4Mux_h
    port map (
            O => \N__30281\,
            I => \N__30273\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__30278\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__5248\ : Odrv4
    port map (
            O => \N__30273\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__5247\ : InMux
    port map (
            O => \N__30268\,
            I => \N__30265\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__30265\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__5245\ : InMux
    port map (
            O => \N__30262\,
            I => \N__30258\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__30261\,
            I => \N__30254\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__30258\,
            I => \N__30251\
        );

    \I__5242\ : InMux
    port map (
            O => \N__30257\,
            I => \N__30248\
        );

    \I__5241\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30245\
        );

    \I__5240\ : Span4Mux_h
    port map (
            O => \N__30251\,
            I => \N__30242\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__30248\,
            I => \current_shift_inst.N_1474_i\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__30245\,
            I => \current_shift_inst.N_1474_i\
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__30242\,
            I => \current_shift_inst.N_1474_i\
        );

    \I__5236\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30232\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__30232\,
            I => \N__30229\
        );

    \I__5234\ : Odrv4
    port map (
            O => \N__30229\,
            I => \current_shift_inst.control_input_18\
        );

    \I__5233\ : InMux
    port map (
            O => \N__30226\,
            I => \N__30223\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__30223\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__5231\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30217\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__30217\,
            I => \N__30214\
        );

    \I__5229\ : Odrv4
    port map (
            O => \N__30214\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__5228\ : InMux
    port map (
            O => \N__30211\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__5227\ : InMux
    port map (
            O => \N__30208\,
            I => \N__30205\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__30205\,
            I => \N__30202\
        );

    \I__5225\ : Odrv4
    port map (
            O => \N__30202\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__5224\ : InMux
    port map (
            O => \N__30199\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__5223\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__30193\,
            I => \N__30190\
        );

    \I__5221\ : Odrv4
    port map (
            O => \N__30190\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__5220\ : InMux
    port map (
            O => \N__30187\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__5219\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30181\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__30181\,
            I => \N__30178\
        );

    \I__5217\ : Odrv4
    port map (
            O => \N__30178\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__5216\ : InMux
    port map (
            O => \N__30175\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__5215\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30169\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__30169\,
            I => \N__30166\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__30166\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__5212\ : InMux
    port map (
            O => \N__30163\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__5211\ : InMux
    port map (
            O => \N__30160\,
            I => \N__30157\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__30154\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__5208\ : InMux
    port map (
            O => \N__30151\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__5207\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30143\
        );

    \I__5206\ : InMux
    port map (
            O => \N__30147\,
            I => \N__30140\
        );

    \I__5205\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30137\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__30143\,
            I => \N__30134\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__30140\,
            I => \N__30129\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__30137\,
            I => \N__30129\
        );

    \I__5201\ : Odrv12
    port map (
            O => \N__30134\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__5200\ : Odrv12
    port map (
            O => \N__30129\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__5199\ : InMux
    port map (
            O => \N__30124\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__5198\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30116\
        );

    \I__5197\ : InMux
    port map (
            O => \N__30120\,
            I => \N__30113\
        );

    \I__5196\ : InMux
    port map (
            O => \N__30119\,
            I => \N__30110\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__30116\,
            I => \N__30105\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__30113\,
            I => \N__30105\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__30110\,
            I => \N__30102\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__30105\,
            I => \N__30099\
        );

    \I__5191\ : Odrv12
    port map (
            O => \N__30102\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__30099\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__5189\ : InMux
    port map (
            O => \N__30094\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__30091\,
            I => \N__30087\
        );

    \I__5187\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30083\
        );

    \I__5186\ : InMux
    port map (
            O => \N__30087\,
            I => \N__30080\
        );

    \I__5185\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30077\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__30083\,
            I => \N__30074\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__30080\,
            I => \N__30069\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__30077\,
            I => \N__30069\
        );

    \I__5181\ : Odrv4
    port map (
            O => \N__30074\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5180\ : Odrv12
    port map (
            O => \N__30069\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__5179\ : InMux
    port map (
            O => \N__30064\,
            I => \bfn_12_10_0_\
        );

    \I__5178\ : InMux
    port map (
            O => \N__30061\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__5177\ : InMux
    port map (
            O => \N__30058\,
            I => \N__30053\
        );

    \I__5176\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30048\
        );

    \I__5175\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30048\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__30053\,
            I => \N__30045\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__30048\,
            I => \N__30042\
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__30045\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__5171\ : Odrv12
    port map (
            O => \N__30042\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__5170\ : InMux
    port map (
            O => \N__30037\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__5169\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30029\
        );

    \I__5168\ : InMux
    port map (
            O => \N__30033\,
            I => \N__30024\
        );

    \I__5167\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30024\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__30029\,
            I => \N__30021\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__30024\,
            I => \N__30018\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__30021\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5163\ : Odrv12
    port map (
            O => \N__30018\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__5162\ : InMux
    port map (
            O => \N__30013\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__5161\ : InMux
    port map (
            O => \N__30010\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__5160\ : InMux
    port map (
            O => \N__30007\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__5159\ : InMux
    port map (
            O => \N__30004\,
            I => \N__30000\
        );

    \I__5158\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29994\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__30000\,
            I => \N__29991\
        );

    \I__5156\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29988\
        );

    \I__5155\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29985\
        );

    \I__5154\ : InMux
    port map (
            O => \N__29997\,
            I => \N__29982\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__29994\,
            I => \N__29979\
        );

    \I__5152\ : Span4Mux_v
    port map (
            O => \N__29991\,
            I => \N__29974\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__29988\,
            I => \N__29974\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__29985\,
            I => \N__29971\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__29982\,
            I => \N__29968\
        );

    \I__5148\ : Span4Mux_h
    port map (
            O => \N__29979\,
            I => \N__29963\
        );

    \I__5147\ : Span4Mux_h
    port map (
            O => \N__29974\,
            I => \N__29963\
        );

    \I__5146\ : Odrv12
    port map (
            O => \N__29971\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5145\ : Odrv4
    port map (
            O => \N__29968\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__29963\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__29956\,
            I => \N__29953\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29953\,
            I => \N__29950\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29950\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0\
        );

    \I__5140\ : CascadeMux
    port map (
            O => \N__29947\,
            I => \N__29944\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29941\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__29941\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29938\,
            I => \N__29935\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__29935\,
            I => \current_shift_inst.PI_CTRL.integrator_i_20\
        );

    \I__5135\ : InMux
    port map (
            O => \N__29932\,
            I => \N__29929\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__29929\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__5133\ : InMux
    port map (
            O => \N__29926\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__5132\ : InMux
    port map (
            O => \N__29923\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__5131\ : InMux
    port map (
            O => \N__29920\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__29917\,
            I => \N__29913\
        );

    \I__5129\ : InMux
    port map (
            O => \N__29916\,
            I => \N__29909\
        );

    \I__5128\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29906\
        );

    \I__5127\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29903\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__29909\,
            I => \N__29900\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29906\,
            I => \N__29895\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__29903\,
            I => \N__29895\
        );

    \I__5123\ : Odrv12
    port map (
            O => \N__29900\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__5122\ : Odrv12
    port map (
            O => \N__29895\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29890\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__29887\,
            I => \N__29883\
        );

    \I__5119\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29879\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29876\
        );

    \I__5117\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29873\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__29879\,
            I => \N__29870\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29865\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__29873\,
            I => \N__29865\
        );

    \I__5113\ : Odrv12
    port map (
            O => \N__29870\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__5112\ : Odrv12
    port map (
            O => \N__29865\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29860\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__29857\,
            I => \N__29853\
        );

    \I__5109\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29849\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29853\,
            I => \N__29846\
        );

    \I__5107\ : CascadeMux
    port map (
            O => \N__29852\,
            I => \N__29843\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__29849\,
            I => \N__29838\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__29846\,
            I => \N__29835\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29832\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__29842\,
            I => \N__29829\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29841\,
            I => \N__29826\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__29838\,
            I => \N__29821\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__29835\,
            I => \N__29821\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29818\
        );

    \I__5098\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29815\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__29826\,
            I => \N__29812\
        );

    \I__5096\ : Odrv4
    port map (
            O => \N__29821\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5095\ : Odrv12
    port map (
            O => \N__29818\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__29815\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__29812\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5092\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29800\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__29800\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0\
        );

    \I__5090\ : CascadeMux
    port map (
            O => \N__29797\,
            I => \N__29794\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29790\
        );

    \I__5088\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29786\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__29790\,
            I => \N__29781\
        );

    \I__5086\ : InMux
    port map (
            O => \N__29789\,
            I => \N__29778\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__29786\,
            I => \N__29775\
        );

    \I__5084\ : InMux
    port map (
            O => \N__29785\,
            I => \N__29770\
        );

    \I__5083\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29770\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__29781\,
            I => \N__29767\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__29778\,
            I => \N__29760\
        );

    \I__5080\ : Span4Mux_h
    port map (
            O => \N__29775\,
            I => \N__29760\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__29770\,
            I => \N__29760\
        );

    \I__5078\ : Odrv4
    port map (
            O => \N__29767\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__29760\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__29755\,
            I => \N__29752\
        );

    \I__5075\ : InMux
    port map (
            O => \N__29752\,
            I => \N__29749\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__29749\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__29746\,
            I => \N__29743\
        );

    \I__5072\ : InMux
    port map (
            O => \N__29743\,
            I => \N__29740\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__29740\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__29737\,
            I => \N__29734\
        );

    \I__5069\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29731\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__29731\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0\
        );

    \I__5067\ : CascadeMux
    port map (
            O => \N__29728\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25_cascade_\
        );

    \I__5066\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29722\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__29722\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0\
        );

    \I__5064\ : InMux
    port map (
            O => \N__29719\,
            I => \N__29715\
        );

    \I__5063\ : InMux
    port map (
            O => \N__29718\,
            I => \N__29711\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29708\
        );

    \I__5061\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29705\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__29711\,
            I => \N__29700\
        );

    \I__5059\ : Span4Mux_h
    port map (
            O => \N__29708\,
            I => \N__29695\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29695\
        );

    \I__5057\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29692\
        );

    \I__5056\ : InMux
    port map (
            O => \N__29703\,
            I => \N__29689\
        );

    \I__5055\ : Span4Mux_h
    port map (
            O => \N__29700\,
            I => \N__29682\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__29695\,
            I => \N__29682\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__29692\,
            I => \N__29682\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__29689\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__29682\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__29677\,
            I => \N__29674\
        );

    \I__5049\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29671\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__29671\,
            I => \N__29668\
        );

    \I__5047\ : Odrv4
    port map (
            O => \N__29668\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0\
        );

    \I__5046\ : CascadeMux
    port map (
            O => \N__29665\,
            I => \N__29662\
        );

    \I__5045\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29659\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__29659\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__29656\,
            I => \N__29653\
        );

    \I__5042\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29649\
        );

    \I__5041\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29646\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__29649\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_14\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__29646\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_14\
        );

    \I__5038\ : CascadeMux
    port map (
            O => \N__29641\,
            I => \N__29638\
        );

    \I__5037\ : InMux
    port map (
            O => \N__29638\,
            I => \N__29634\
        );

    \I__5036\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29630\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__29634\,
            I => \N__29627\
        );

    \I__5034\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29624\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__29630\,
            I => \N__29620\
        );

    \I__5032\ : Span4Mux_v
    port map (
            O => \N__29627\,
            I => \N__29615\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__29624\,
            I => \N__29615\
        );

    \I__5030\ : InMux
    port map (
            O => \N__29623\,
            I => \N__29611\
        );

    \I__5029\ : Span4Mux_h
    port map (
            O => \N__29620\,
            I => \N__29608\
        );

    \I__5028\ : Span4Mux_h
    port map (
            O => \N__29615\,
            I => \N__29605\
        );

    \I__5027\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29602\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__29611\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__29608\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__29605\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__29602\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29593\,
            I => \N__29590\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__29590\,
            I => \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9\
        );

    \I__5020\ : CascadeMux
    port map (
            O => \N__29587\,
            I => \N__29584\
        );

    \I__5019\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29579\
        );

    \I__5018\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29576\
        );

    \I__5017\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29573\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__29579\,
            I => \N__29570\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__29576\,
            I => \N__29567\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__29573\,
            I => \N__29563\
        );

    \I__5013\ : Span4Mux_v
    port map (
            O => \N__29570\,
            I => \N__29560\
        );

    \I__5012\ : Span4Mux_h
    port map (
            O => \N__29567\,
            I => \N__29556\
        );

    \I__5011\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29553\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__29563\,
            I => \N__29550\
        );

    \I__5009\ : Span4Mux_h
    port map (
            O => \N__29560\,
            I => \N__29547\
        );

    \I__5008\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29544\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__29556\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__29553\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__29550\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__29547\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__29544\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__5002\ : CascadeMux
    port map (
            O => \N__29533\,
            I => \N__29530\
        );

    \I__5001\ : InMux
    port map (
            O => \N__29530\,
            I => \N__29527\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__29527\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8\
        );

    \I__4999\ : CascadeMux
    port map (
            O => \N__29524\,
            I => \N__29521\
        );

    \I__4998\ : InMux
    port map (
            O => \N__29521\,
            I => \N__29518\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__29518\,
            I => \N__29515\
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__29515\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0\
        );

    \I__4995\ : CascadeMux
    port map (
            O => \N__29512\,
            I => \N__29509\
        );

    \I__4994\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29506\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__29506\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0\
        );

    \I__4992\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29500\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__29500\,
            I => \current_shift_inst.PI_CTRL.integrator_i_10\
        );

    \I__4990\ : InMux
    port map (
            O => \N__29497\,
            I => \N__29494\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__29494\,
            I => \current_shift_inst.PI_CTRL.integrator_i_13\
        );

    \I__4988\ : InMux
    port map (
            O => \N__29491\,
            I => \N__29487\
        );

    \I__4987\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29484\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__29487\,
            I => \N__29478\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29475\
        );

    \I__4984\ : CascadeMux
    port map (
            O => \N__29483\,
            I => \N__29472\
        );

    \I__4983\ : CascadeMux
    port map (
            O => \N__29482\,
            I => \N__29469\
        );

    \I__4982\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29466\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__29478\,
            I => \N__29463\
        );

    \I__4980\ : Span4Mux_h
    port map (
            O => \N__29475\,
            I => \N__29460\
        );

    \I__4979\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29455\
        );

    \I__4978\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29455\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__29466\,
            I => \N__29452\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__29463\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4975\ : Odrv4
    port map (
            O => \N__29460\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__29455\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4973\ : Odrv4
    port map (
            O => \N__29452\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4972\ : CascadeMux
    port map (
            O => \N__29443\,
            I => \N__29440\
        );

    \I__4971\ : InMux
    port map (
            O => \N__29440\,
            I => \N__29437\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__29437\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0\
        );

    \I__4969\ : CascadeMux
    port map (
            O => \N__29434\,
            I => \N__29431\
        );

    \I__4968\ : InMux
    port map (
            O => \N__29431\,
            I => \N__29427\
        );

    \I__4967\ : InMux
    port map (
            O => \N__29430\,
            I => \N__29424\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__29427\,
            I => \N__29421\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__29424\,
            I => \N__29417\
        );

    \I__4964\ : Span4Mux_v
    port map (
            O => \N__29421\,
            I => \N__29413\
        );

    \I__4963\ : InMux
    port map (
            O => \N__29420\,
            I => \N__29410\
        );

    \I__4962\ : Span4Mux_v
    port map (
            O => \N__29417\,
            I => \N__29407\
        );

    \I__4961\ : InMux
    port map (
            O => \N__29416\,
            I => \N__29404\
        );

    \I__4960\ : Span4Mux_h
    port map (
            O => \N__29413\,
            I => \N__29401\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__29410\,
            I => \N__29398\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__29407\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__29404\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__29401\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__29398\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__29389\,
            I => \N__29386\
        );

    \I__4953\ : InMux
    port map (
            O => \N__29386\,
            I => \N__29383\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__29383\,
            I => \N__29380\
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__29380\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5\
        );

    \I__4950\ : InMux
    port map (
            O => \N__29377\,
            I => \N__29374\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29374\,
            I => \N__29370\
        );

    \I__4948\ : InMux
    port map (
            O => \N__29373\,
            I => \N__29367\
        );

    \I__4947\ : Span4Mux_v
    port map (
            O => \N__29370\,
            I => \N__29364\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__29367\,
            I => \N__29361\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__29364\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__4944\ : Odrv12
    port map (
            O => \N__29361\,
            I => \current_shift_inst.PI_CTRL.integrator_i_0\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__29356\,
            I => \N__29353\
        );

    \I__4942\ : InMux
    port map (
            O => \N__29353\,
            I => \N__29350\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__29350\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4\
        );

    \I__4940\ : CascadeMux
    port map (
            O => \N__29347\,
            I => \N__29343\
        );

    \I__4939\ : CascadeMux
    port map (
            O => \N__29346\,
            I => \N__29340\
        );

    \I__4938\ : InMux
    port map (
            O => \N__29343\,
            I => \N__29335\
        );

    \I__4937\ : InMux
    port map (
            O => \N__29340\,
            I => \N__29332\
        );

    \I__4936\ : InMux
    port map (
            O => \N__29339\,
            I => \N__29329\
        );

    \I__4935\ : InMux
    port map (
            O => \N__29338\,
            I => \N__29325\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__29335\,
            I => \N__29322\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__29332\,
            I => \N__29319\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__29329\,
            I => \N__29316\
        );

    \I__4931\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29313\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__29325\,
            I => \N__29310\
        );

    \I__4929\ : Span4Mux_h
    port map (
            O => \N__29322\,
            I => \N__29307\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__29319\,
            I => \N__29304\
        );

    \I__4927\ : Span4Mux_h
    port map (
            O => \N__29316\,
            I => \N__29297\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__29313\,
            I => \N__29297\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__29310\,
            I => \N__29297\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__29307\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__29304\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__29297\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__29290\,
            I => \N__29287\
        );

    \I__4920\ : InMux
    port map (
            O => \N__29287\,
            I => \N__29284\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__29284\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10\
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__29281\,
            I => \N__29278\
        );

    \I__4917\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29275\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__29275\,
            I => \N__29272\
        );

    \I__4915\ : Span4Mux_h
    port map (
            O => \N__29272\,
            I => \N__29269\
        );

    \I__4914\ : Odrv4
    port map (
            O => \N__29269\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13\
        );

    \I__4913\ : InMux
    port map (
            O => \N__29266\,
            I => \N__29263\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__29263\,
            I => \N__29258\
        );

    \I__4911\ : InMux
    port map (
            O => \N__29262\,
            I => \N__29254\
        );

    \I__4910\ : InMux
    port map (
            O => \N__29261\,
            I => \N__29251\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__29258\,
            I => \N__29248\
        );

    \I__4908\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29245\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__29254\,
            I => \N__29242\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29239\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__29248\,
            I => \N__29234\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__29245\,
            I => \N__29234\
        );

    \I__4903\ : Span4Mux_v
    port map (
            O => \N__29242\,
            I => \N__29229\
        );

    \I__4902\ : Span4Mux_h
    port map (
            O => \N__29239\,
            I => \N__29229\
        );

    \I__4901\ : Odrv4
    port map (
            O => \N__29234\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__29229\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__4899\ : CascadeMux
    port map (
            O => \N__29224\,
            I => \N__29221\
        );

    \I__4898\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29218\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__29218\,
            I => \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6\
        );

    \I__4896\ : CascadeMux
    port map (
            O => \N__29215\,
            I => \N__29211\
        );

    \I__4895\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29208\
        );

    \I__4894\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29205\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__29208\,
            I => \N__29200\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__29205\,
            I => \N__29197\
        );

    \I__4891\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29194\
        );

    \I__4890\ : InMux
    port map (
            O => \N__29203\,
            I => \N__29190\
        );

    \I__4889\ : Span4Mux_v
    port map (
            O => \N__29200\,
            I => \N__29183\
        );

    \I__4888\ : Span4Mux_v
    port map (
            O => \N__29197\,
            I => \N__29183\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__29194\,
            I => \N__29183\
        );

    \I__4886\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29180\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__29190\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__29183\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__29180\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4882\ : CascadeMux
    port map (
            O => \N__29173\,
            I => \N__29170\
        );

    \I__4881\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29167\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__29167\,
            I => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0\
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__29164\,
            I => \N__29161\
        );

    \I__4878\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29158\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__29158\,
            I => \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11\
        );

    \I__4876\ : InMux
    port map (
            O => \N__29155\,
            I => \N__29151\
        );

    \I__4875\ : InMux
    port map (
            O => \N__29154\,
            I => \N__29148\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__29151\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__29148\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__4872\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29139\
        );

    \I__4871\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29136\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__29139\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__29136\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__4868\ : InMux
    port map (
            O => \N__29131\,
            I => \N__29128\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__29128\,
            I => \N__29125\
        );

    \I__4866\ : Odrv12
    port map (
            O => \N__29125\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df28\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__29122\,
            I => \N__29119\
        );

    \I__4864\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29116\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__29116\,
            I => \N__29110\
        );

    \I__4862\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29107\
        );

    \I__4861\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29104\
        );

    \I__4860\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29101\
        );

    \I__4859\ : Span4Mux_h
    port map (
            O => \N__29110\,
            I => \N__29096\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__29107\,
            I => \N__29096\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__29104\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__29101\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__29096\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__4854\ : InMux
    port map (
            O => \N__29089\,
            I => \N__29084\
        );

    \I__4853\ : InMux
    port map (
            O => \N__29088\,
            I => \N__29081\
        );

    \I__4852\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29078\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__29084\,
            I => \N__29075\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__29081\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__29078\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__29075\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__4847\ : InMux
    port map (
            O => \N__29068\,
            I => \N__29065\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N__29062\
        );

    \I__4845\ : Odrv4
    port map (
            O => \N__29062\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__4844\ : InMux
    port map (
            O => \N__29059\,
            I => \N__29056\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__29056\,
            I => \N__29052\
        );

    \I__4842\ : InMux
    port map (
            O => \N__29055\,
            I => \N__29049\
        );

    \I__4841\ : Span12Mux_v
    port map (
            O => \N__29052\,
            I => \N__29044\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__29041\
        );

    \I__4839\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29038\
        );

    \I__4838\ : InMux
    port map (
            O => \N__29047\,
            I => \N__29035\
        );

    \I__4837\ : Span12Mux_v
    port map (
            O => \N__29044\,
            I => \N__29032\
        );

    \I__4836\ : Span12Mux_v
    port map (
            O => \N__29041\,
            I => \N__29029\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__29038\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__29035\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__4833\ : Odrv12
    port map (
            O => \N__29032\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__4832\ : Odrv12
    port map (
            O => \N__29029\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__4831\ : ClkMux
    port map (
            O => \N__29020\,
            I => \N__29014\
        );

    \I__4830\ : ClkMux
    port map (
            O => \N__29019\,
            I => \N__29014\
        );

    \I__4829\ : GlobalMux
    port map (
            O => \N__29014\,
            I => \N__29011\
        );

    \I__4828\ : gio2CtrlBuf
    port map (
            O => \N__29011\,
            I => delay_tr_input_c_g
        );

    \I__4827\ : InMux
    port map (
            O => \N__29008\,
            I => \N__29005\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__29005\,
            I => \N__29002\
        );

    \I__4825\ : Span4Mux_v
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__4824\ : Span4Mux_v
    port map (
            O => \N__28999\,
            I => \N__28994\
        );

    \I__4823\ : InMux
    port map (
            O => \N__28998\,
            I => \N__28991\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28988\
        );

    \I__4821\ : Span4Mux_v
    port map (
            O => \N__28994\,
            I => \N__28985\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__28991\,
            I => \N__28982\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28979\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__28985\,
            I => \N__28976\
        );

    \I__4817\ : Sp12to4
    port map (
            O => \N__28982\,
            I => \N__28973\
        );

    \I__4816\ : Span12Mux_v
    port map (
            O => \N__28979\,
            I => \N__28970\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__28976\,
            I => \N__28967\
        );

    \I__4814\ : Odrv12
    port map (
            O => \N__28973\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__4813\ : Odrv12
    port map (
            O => \N__28970\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__28967\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__4811\ : IoInMux
    port map (
            O => \N__28960\,
            I => \N__28957\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__28957\,
            I => \N__28954\
        );

    \I__4809\ : Odrv4
    port map (
            O => \N__28954\,
            I => \delay_measurement_inst.delay_tr_timer.N_399_i\
        );

    \I__4808\ : CascadeMux
    port map (
            O => \N__28951\,
            I => \N__28948\
        );

    \I__4807\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28945\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__28945\,
            I => \N__28942\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__28942\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__4804\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28933\
        );

    \I__4803\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28933\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__28933\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__28930\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28924\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__28924\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__4798\ : InMux
    port map (
            O => \N__28921\,
            I => \N__28909\
        );

    \I__4797\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28909\
        );

    \I__4796\ : InMux
    port map (
            O => \N__28919\,
            I => \N__28909\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28918\,
            I => \N__28909\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__28909\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__28906\,
            I => \N__28902\
        );

    \I__4792\ : CascadeMux
    port map (
            O => \N__28905\,
            I => \N__28899\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28894\
        );

    \I__4790\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28894\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__28894\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__4788\ : InMux
    port map (
            O => \N__28891\,
            I => \N__28888\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__28888\,
            I => \N__28885\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__28885\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__4785\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28878\
        );

    \I__4784\ : InMux
    port map (
            O => \N__28881\,
            I => \N__28875\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__28878\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__28875\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__4781\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28866\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28869\,
            I => \N__28863\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__28866\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__28863\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__4777\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28855\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__28855\,
            I => \N__28852\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__28852\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df20\
        );

    \I__4774\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28845\
        );

    \I__4773\ : InMux
    port map (
            O => \N__28848\,
            I => \N__28842\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__28845\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__28842\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28837\,
            I => \N__28833\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28836\,
            I => \N__28830\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__28833\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__28830\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__4766\ : InMux
    port map (
            O => \N__28825\,
            I => \N__28822\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__28822\,
            I => \N__28819\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__28819\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df22\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28812\
        );

    \I__4762\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28809\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__28812\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__28809\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__4759\ : InMux
    port map (
            O => \N__28804\,
            I => \N__28800\
        );

    \I__4758\ : InMux
    port map (
            O => \N__28803\,
            I => \N__28797\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__28800\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__28797\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__4755\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28789\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__28789\,
            I => \N__28786\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__28786\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df24\
        );

    \I__4752\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28779\
        );

    \I__4751\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28776\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__28779\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__28776\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__4748\ : InMux
    port map (
            O => \N__28771\,
            I => \N__28767\
        );

    \I__4747\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28764\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__28767\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28764\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__4744\ : InMux
    port map (
            O => \N__28759\,
            I => \N__28756\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__28756\,
            I => \N__28753\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__28753\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df26\
        );

    \I__4741\ : InMux
    port map (
            O => \N__28750\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28\
        );

    \I__4740\ : InMux
    port map (
            O => \N__28747\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__28744\,
            I => \N__28741\
        );

    \I__4738\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28738\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__28738\,
            I => \N__28735\
        );

    \I__4736\ : Odrv4
    port map (
            O => \N__28735\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28\
        );

    \I__4735\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28726\
        );

    \I__4734\ : InMux
    port map (
            O => \N__28731\,
            I => \N__28726\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__28726\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__28723\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__28720\,
            I => \N__28715\
        );

    \I__4730\ : InMux
    port map (
            O => \N__28719\,
            I => \N__28712\
        );

    \I__4729\ : InMux
    port map (
            O => \N__28718\,
            I => \N__28709\
        );

    \I__4728\ : InMux
    port map (
            O => \N__28715\,
            I => \N__28706\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__28712\,
            I => \N__28703\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__28709\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__28706\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4724\ : Odrv4
    port map (
            O => \N__28703\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4723\ : InMux
    port map (
            O => \N__28696\,
            I => \N__28692\
        );

    \I__4722\ : InMux
    port map (
            O => \N__28695\,
            I => \N__28689\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__28692\,
            I => \N__28686\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__28689\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__28686\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4718\ : CascadeMux
    port map (
            O => \N__28681\,
            I => \N__28678\
        );

    \I__4717\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28675\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__28675\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__4715\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28668\
        );

    \I__4714\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28665\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__28668\,
            I => \N__28662\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__28665\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__28662\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4710\ : CascadeMux
    port map (
            O => \N__28657\,
            I => \N__28654\
        );

    \I__4709\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28651\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__28651\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__4707\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28644\
        );

    \I__4706\ : InMux
    port map (
            O => \N__28647\,
            I => \N__28641\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__28644\,
            I => \N__28638\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__28641\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__28638\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4702\ : CascadeMux
    port map (
            O => \N__28633\,
            I => \N__28630\
        );

    \I__4701\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28627\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__28627\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__4699\ : InMux
    port map (
            O => \N__28624\,
            I => \N__28620\
        );

    \I__4698\ : InMux
    port map (
            O => \N__28623\,
            I => \N__28617\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__28620\,
            I => \N__28614\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__28617\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__28614\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__28609\,
            I => \N__28606\
        );

    \I__4693\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28603\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__28603\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__4691\ : InMux
    port map (
            O => \N__28600\,
            I => \N__28596\
        );

    \I__4690\ : InMux
    port map (
            O => \N__28599\,
            I => \N__28593\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__28596\,
            I => \N__28590\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__28593\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4687\ : Odrv4
    port map (
            O => \N__28590\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4686\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28582\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__28582\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__4684\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28575\
        );

    \I__4683\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28572\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__28575\,
            I => \N__28569\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__28572\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__28569\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__28564\,
            I => \N__28561\
        );

    \I__4678\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28558\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__28558\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__4676\ : InMux
    port map (
            O => \N__28555\,
            I => \N__28551\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28548\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__28551\,
            I => \N__28545\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__28548\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__28545\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4671\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28537\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__28537\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__4669\ : InMux
    port map (
            O => \N__28534\,
            I => \N__28530\
        );

    \I__4668\ : InMux
    port map (
            O => \N__28533\,
            I => \N__28527\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__28530\,
            I => \N__28524\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__28527\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__28524\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__28519\,
            I => \N__28516\
        );

    \I__4663\ : InMux
    port map (
            O => \N__28516\,
            I => \N__28513\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__28513\,
            I => \N__28510\
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__28510\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__4660\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28503\
        );

    \I__4659\ : InMux
    port map (
            O => \N__28506\,
            I => \N__28500\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__28503\,
            I => \N__28497\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__28500\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__28497\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__28492\,
            I => \N__28489\
        );

    \I__4654\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28486\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__28486\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__4652\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28479\
        );

    \I__4651\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28476\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__28479\,
            I => \N__28473\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__28476\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__28473\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4647\ : InMux
    port map (
            O => \N__28468\,
            I => \N__28465\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__28465\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__4645\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28458\
        );

    \I__4644\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28455\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__28458\,
            I => \N__28452\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__28455\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__28452\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4640\ : CascadeMux
    port map (
            O => \N__28447\,
            I => \N__28444\
        );

    \I__4639\ : InMux
    port map (
            O => \N__28444\,
            I => \N__28441\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__28441\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__4637\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28435\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__28435\,
            I => \N__28431\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28434\,
            I => \N__28428\
        );

    \I__4634\ : Span4Mux_h
    port map (
            O => \N__28431\,
            I => \N__28425\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__28428\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4632\ : Odrv4
    port map (
            O => \N__28425\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4631\ : CascadeMux
    port map (
            O => \N__28420\,
            I => \N__28417\
        );

    \I__4630\ : InMux
    port map (
            O => \N__28417\,
            I => \N__28414\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__28414\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__4628\ : InMux
    port map (
            O => \N__28411\,
            I => \N__28407\
        );

    \I__4627\ : InMux
    port map (
            O => \N__28410\,
            I => \N__28404\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__28407\,
            I => \N__28401\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__28404\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4624\ : Odrv4
    port map (
            O => \N__28401\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4623\ : CascadeMux
    port map (
            O => \N__28396\,
            I => \N__28393\
        );

    \I__4622\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28390\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__28390\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__28387\,
            I => \N__28384\
        );

    \I__4619\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28381\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__28381\,
            I => \N__28378\
        );

    \I__4617\ : Span4Mux_h
    port map (
            O => \N__28378\,
            I => \N__28375\
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__28375\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__4615\ : InMux
    port map (
            O => \N__28372\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__4614\ : InMux
    port map (
            O => \N__28369\,
            I => \N__28366\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__28366\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__4612\ : InMux
    port map (
            O => \N__28363\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__4611\ : CascadeMux
    port map (
            O => \N__28360\,
            I => \N__28357\
        );

    \I__4610\ : InMux
    port map (
            O => \N__28357\,
            I => \N__28354\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__28354\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__4608\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28348\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__28348\,
            I => \N__28345\
        );

    \I__4606\ : Odrv12
    port map (
            O => \N__28345\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__4605\ : InMux
    port map (
            O => \N__28342\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__4604\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28336\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__28336\,
            I => \N__28333\
        );

    \I__4602\ : Span4Mux_v
    port map (
            O => \N__28333\,
            I => \N__28330\
        );

    \I__4601\ : Odrv4
    port map (
            O => \N__28330\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__4600\ : InMux
    port map (
            O => \N__28327\,
            I => \N__28324\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__28324\,
            I => \N__28321\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__28321\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__4597\ : InMux
    port map (
            O => \N__28318\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__4596\ : InMux
    port map (
            O => \N__28315\,
            I => \N__28305\
        );

    \I__4595\ : InMux
    port map (
            O => \N__28314\,
            I => \N__28297\
        );

    \I__4594\ : InMux
    port map (
            O => \N__28313\,
            I => \N__28290\
        );

    \I__4593\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28290\
        );

    \I__4592\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28290\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__28310\,
            I => \N__28278\
        );

    \I__4590\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28263\
        );

    \I__4589\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28260\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__28305\,
            I => \N__28257\
        );

    \I__4587\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28254\
        );

    \I__4586\ : InMux
    port map (
            O => \N__28303\,
            I => \N__28245\
        );

    \I__4585\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28245\
        );

    \I__4584\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28245\
        );

    \I__4583\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28245\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28240\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__28290\,
            I => \N__28240\
        );

    \I__4580\ : InMux
    port map (
            O => \N__28289\,
            I => \N__28237\
        );

    \I__4579\ : InMux
    port map (
            O => \N__28288\,
            I => \N__28230\
        );

    \I__4578\ : InMux
    port map (
            O => \N__28287\,
            I => \N__28230\
        );

    \I__4577\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28230\
        );

    \I__4576\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28221\
        );

    \I__4575\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28221\
        );

    \I__4574\ : InMux
    port map (
            O => \N__28283\,
            I => \N__28221\
        );

    \I__4573\ : InMux
    port map (
            O => \N__28282\,
            I => \N__28221\
        );

    \I__4572\ : InMux
    port map (
            O => \N__28281\,
            I => \N__28213\
        );

    \I__4571\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28213\
        );

    \I__4570\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28213\
        );

    \I__4569\ : CascadeMux
    port map (
            O => \N__28276\,
            I => \N__28208\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__28275\,
            I => \N__28204\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__28274\,
            I => \N__28200\
        );

    \I__4566\ : CascadeMux
    port map (
            O => \N__28273\,
            I => \N__28196\
        );

    \I__4565\ : CascadeMux
    port map (
            O => \N__28272\,
            I => \N__28192\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__28271\,
            I => \N__28188\
        );

    \I__4563\ : CascadeMux
    port map (
            O => \N__28270\,
            I => \N__28184\
        );

    \I__4562\ : CascadeMux
    port map (
            O => \N__28269\,
            I => \N__28180\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__28268\,
            I => \N__28176\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__28267\,
            I => \N__28172\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__28266\,
            I => \N__28168\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__28263\,
            I => \N__28161\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__28260\,
            I => \N__28158\
        );

    \I__4556\ : Span4Mux_s1_v
    port map (
            O => \N__28257\,
            I => \N__28153\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__28254\,
            I => \N__28153\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__28245\,
            I => \N__28150\
        );

    \I__4553\ : Span4Mux_v
    port map (
            O => \N__28240\,
            I => \N__28141\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__28237\,
            I => \N__28141\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__28230\,
            I => \N__28141\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__28221\,
            I => \N__28141\
        );

    \I__4549\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28138\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__28213\,
            I => \N__28135\
        );

    \I__4547\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28132\
        );

    \I__4546\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28117\
        );

    \I__4545\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28117\
        );

    \I__4544\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28117\
        );

    \I__4543\ : InMux
    port map (
            O => \N__28204\,
            I => \N__28117\
        );

    \I__4542\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28117\
        );

    \I__4541\ : InMux
    port map (
            O => \N__28200\,
            I => \N__28117\
        );

    \I__4540\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28117\
        );

    \I__4539\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28100\
        );

    \I__4538\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28100\
        );

    \I__4537\ : InMux
    port map (
            O => \N__28192\,
            I => \N__28100\
        );

    \I__4536\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28100\
        );

    \I__4535\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28100\
        );

    \I__4534\ : InMux
    port map (
            O => \N__28187\,
            I => \N__28100\
        );

    \I__4533\ : InMux
    port map (
            O => \N__28184\,
            I => \N__28100\
        );

    \I__4532\ : InMux
    port map (
            O => \N__28183\,
            I => \N__28100\
        );

    \I__4531\ : InMux
    port map (
            O => \N__28180\,
            I => \N__28083\
        );

    \I__4530\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28083\
        );

    \I__4529\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28083\
        );

    \I__4528\ : InMux
    port map (
            O => \N__28175\,
            I => \N__28083\
        );

    \I__4527\ : InMux
    port map (
            O => \N__28172\,
            I => \N__28083\
        );

    \I__4526\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28083\
        );

    \I__4525\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28083\
        );

    \I__4524\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28083\
        );

    \I__4523\ : CascadeMux
    port map (
            O => \N__28166\,
            I => \N__28079\
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__28165\,
            I => \N__28075\
        );

    \I__4521\ : CascadeMux
    port map (
            O => \N__28164\,
            I => \N__28071\
        );

    \I__4520\ : Span12Mux_v
    port map (
            O => \N__28161\,
            I => \N__28067\
        );

    \I__4519\ : Span12Mux_s1_h
    port map (
            O => \N__28158\,
            I => \N__28062\
        );

    \I__4518\ : Sp12to4
    port map (
            O => \N__28153\,
            I => \N__28062\
        );

    \I__4517\ : Sp12to4
    port map (
            O => \N__28150\,
            I => \N__28057\
        );

    \I__4516\ : Sp12to4
    port map (
            O => \N__28141\,
            I => \N__28057\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__28138\,
            I => \N__28054\
        );

    \I__4514\ : Span4Mux_h
    port map (
            O => \N__28135\,
            I => \N__28051\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__28132\,
            I => \N__28048\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__28117\,
            I => \N__28041\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__28100\,
            I => \N__28041\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__28083\,
            I => \N__28041\
        );

    \I__4509\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28026\
        );

    \I__4508\ : InMux
    port map (
            O => \N__28079\,
            I => \N__28026\
        );

    \I__4507\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28026\
        );

    \I__4506\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28026\
        );

    \I__4505\ : InMux
    port map (
            O => \N__28074\,
            I => \N__28026\
        );

    \I__4504\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28026\
        );

    \I__4503\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28026\
        );

    \I__4502\ : Span12Mux_h
    port map (
            O => \N__28067\,
            I => \N__28019\
        );

    \I__4501\ : Span12Mux_v
    port map (
            O => \N__28062\,
            I => \N__28019\
        );

    \I__4500\ : Span12Mux_v
    port map (
            O => \N__28057\,
            I => \N__28019\
        );

    \I__4499\ : Span4Mux_v
    port map (
            O => \N__28054\,
            I => \N__28016\
        );

    \I__4498\ : Span4Mux_v
    port map (
            O => \N__28051\,
            I => \N__28007\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__28048\,
            I => \N__28007\
        );

    \I__4496\ : Span4Mux_v
    port map (
            O => \N__28041\,
            I => \N__28007\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__28026\,
            I => \N__28007\
        );

    \I__4494\ : Odrv12
    port map (
            O => \N__28019\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__28016\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__28007\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__28000\,
            I => \N__27997\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27992\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__27996\,
            I => \N__27987\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27995\,
            I => \N__27984\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__27992\,
            I => \N__27981\
        );

    \I__4486\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27976\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27990\,
            I => \N__27976\
        );

    \I__4484\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27973\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27969\
        );

    \I__4482\ : Span4Mux_h
    port map (
            O => \N__27981\,
            I => \N__27964\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__27976\,
            I => \N__27964\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__27973\,
            I => \N__27961\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27972\,
            I => \N__27958\
        );

    \I__4478\ : Span4Mux_h
    port map (
            O => \N__27969\,
            I => \N__27955\
        );

    \I__4477\ : Span4Mux_v
    port map (
            O => \N__27964\,
            I => \N__27952\
        );

    \I__4476\ : Odrv4
    port map (
            O => \N__27961\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27958\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__4474\ : Odrv4
    port map (
            O => \N__27955\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__27952\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__4472\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27939\
        );

    \I__4471\ : CascadeMux
    port map (
            O => \N__27942\,
            I => \N__27936\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__27939\,
            I => \N__27933\
        );

    \I__4469\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27930\
        );

    \I__4468\ : Odrv12
    port map (
            O => \N__27933\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__27930\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__4466\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27921\
        );

    \I__4465\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27918\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__27921\,
            I => \N__27915\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__27918\,
            I => \N__27912\
        );

    \I__4462\ : Span4Mux_v
    port map (
            O => \N__27915\,
            I => \N__27907\
        );

    \I__4461\ : Span4Mux_h
    port map (
            O => \N__27912\,
            I => \N__27907\
        );

    \I__4460\ : Odrv4
    port map (
            O => \N__27907\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__27904\,
            I => \N__27901\
        );

    \I__4458\ : InMux
    port map (
            O => \N__27901\,
            I => \N__27898\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__27898\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__4456\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27892\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__27892\,
            I => \N__27888\
        );

    \I__4454\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27885\
        );

    \I__4453\ : Span4Mux_h
    port map (
            O => \N__27888\,
            I => \N__27882\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__27885\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4451\ : Odrv4
    port map (
            O => \N__27882\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4450\ : InMux
    port map (
            O => \N__27877\,
            I => \N__27874\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__27874\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__27871\,
            I => \N__27868\
        );

    \I__4447\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27865\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__27865\,
            I => \N__27862\
        );

    \I__4445\ : Span4Mux_v
    port map (
            O => \N__27862\,
            I => \N__27859\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__27859\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27853\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__27853\,
            I => \N__27850\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__27850\,
            I => \N__27847\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__27847\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__4439\ : InMux
    port map (
            O => \N__27844\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27838\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__27838\,
            I => \N__27835\
        );

    \I__4436\ : Span4Mux_v
    port map (
            O => \N__27835\,
            I => \N__27832\
        );

    \I__4435\ : Odrv4
    port map (
            O => \N__27832\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__4434\ : InMux
    port map (
            O => \N__27829\,
            I => \N__27826\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__27826\,
            I => \N__27823\
        );

    \I__4432\ : Odrv12
    port map (
            O => \N__27823\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27820\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__4430\ : InMux
    port map (
            O => \N__27817\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27814\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__4428\ : InMux
    port map (
            O => \N__27811\,
            I => \bfn_11_18_0_\
        );

    \I__4427\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__27805\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__4425\ : InMux
    port map (
            O => \N__27802\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__27799\,
            I => \N__27796\
        );

    \I__4423\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27793\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__27793\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__4421\ : InMux
    port map (
            O => \N__27790\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27784\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__27784\,
            I => \N__27781\
        );

    \I__4418\ : Odrv12
    port map (
            O => \N__27781\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__4417\ : InMux
    port map (
            O => \N__27778\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__4416\ : InMux
    port map (
            O => \N__27775\,
            I => \N__27772\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__27772\,
            I => \N__27769\
        );

    \I__4414\ : Odrv12
    port map (
            O => \N__27769\,
            I => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__27766\,
            I => \N__27763\
        );

    \I__4412\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27760\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27760\,
            I => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\
        );

    \I__4410\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27754\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__27754\,
            I => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__27751\,
            I => \N__27748\
        );

    \I__4407\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27745\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__27745\,
            I => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\
        );

    \I__4405\ : InMux
    port map (
            O => \N__27742\,
            I => \N__27739\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__27739\,
            I => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\
        );

    \I__4403\ : CascadeMux
    port map (
            O => \N__27736\,
            I => \N__27733\
        );

    \I__4402\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27730\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__27730\,
            I => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\
        );

    \I__4400\ : CascadeMux
    port map (
            O => \N__27727\,
            I => \N__27724\
        );

    \I__4399\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27721\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27721\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__4397\ : CascadeMux
    port map (
            O => \N__27718\,
            I => \N__27715\
        );

    \I__4396\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27712\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__27712\,
            I => \N__27709\
        );

    \I__4394\ : Odrv4
    port map (
            O => \N__27709\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__4393\ : CascadeMux
    port map (
            O => \N__27706\,
            I => \N__27703\
        );

    \I__4392\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27700\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__27700\,
            I => \N__27697\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__27697\,
            I => \N__27694\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__27694\,
            I => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\
        );

    \I__4388\ : InMux
    port map (
            O => \N__27691\,
            I => \N__27688\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__27688\,
            I => \N__27685\
        );

    \I__4386\ : Span4Mux_v
    port map (
            O => \N__27685\,
            I => \N__27682\
        );

    \I__4385\ : Odrv4
    port map (
            O => \N__27682\,
            I => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__27679\,
            I => \N__27676\
        );

    \I__4383\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27673\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__27673\,
            I => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\
        );

    \I__4381\ : InMux
    port map (
            O => \N__27670\,
            I => \N__27667\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__27667\,
            I => \N__27663\
        );

    \I__4379\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27660\
        );

    \I__4378\ : Span4Mux_v
    port map (
            O => \N__27663\,
            I => \N__27654\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__27660\,
            I => \N__27654\
        );

    \I__4376\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27651\
        );

    \I__4375\ : Span4Mux_h
    port map (
            O => \N__27654\,
            I => \N__27648\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__27651\,
            I => \N__27645\
        );

    \I__4373\ : Span4Mux_v
    port map (
            O => \N__27648\,
            I => \N__27642\
        );

    \I__4372\ : Span4Mux_h
    port map (
            O => \N__27645\,
            I => \N__27639\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__27642\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__4370\ : Odrv4
    port map (
            O => \N__27639\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__4369\ : CEMux
    port map (
            O => \N__27634\,
            I => \N__27607\
        );

    \I__4368\ : CEMux
    port map (
            O => \N__27633\,
            I => \N__27607\
        );

    \I__4367\ : CEMux
    port map (
            O => \N__27632\,
            I => \N__27607\
        );

    \I__4366\ : CEMux
    port map (
            O => \N__27631\,
            I => \N__27607\
        );

    \I__4365\ : CEMux
    port map (
            O => \N__27630\,
            I => \N__27607\
        );

    \I__4364\ : CEMux
    port map (
            O => \N__27629\,
            I => \N__27607\
        );

    \I__4363\ : CEMux
    port map (
            O => \N__27628\,
            I => \N__27607\
        );

    \I__4362\ : CEMux
    port map (
            O => \N__27627\,
            I => \N__27607\
        );

    \I__4361\ : CEMux
    port map (
            O => \N__27626\,
            I => \N__27607\
        );

    \I__4360\ : GlobalMux
    port map (
            O => \N__27607\,
            I => \N__27604\
        );

    \I__4359\ : gio2CtrlBuf
    port map (
            O => \N__27604\,
            I => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \I__4358\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27594\
        );

    \I__4357\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27594\
        );

    \I__4356\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27591\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__27594\,
            I => \N__27588\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__27591\,
            I => \N__27585\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__27588\,
            I => \N__27582\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__27585\,
            I => \N__27579\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__27582\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__4350\ : Odrv4
    port map (
            O => \N__27579\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__27574\,
            I => \N__27571\
        );

    \I__4348\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27565\
        );

    \I__4347\ : InMux
    port map (
            O => \N__27570\,
            I => \N__27565\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__27565\,
            I => \N__27562\
        );

    \I__4345\ : Span4Mux_v
    port map (
            O => \N__27562\,
            I => \N__27559\
        );

    \I__4344\ : Span4Mux_h
    port map (
            O => \N__27559\,
            I => \N__27554\
        );

    \I__4343\ : InMux
    port map (
            O => \N__27558\,
            I => \N__27551\
        );

    \I__4342\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27548\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__27554\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__27551\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__27548\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__27541\,
            I => \N__27538\
        );

    \I__4337\ : InMux
    port map (
            O => \N__27538\,
            I => \N__27535\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__27535\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__4335\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27529\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__27529\,
            I => \N__27524\
        );

    \I__4333\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27521\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__27527\,
            I => \N__27518\
        );

    \I__4331\ : Span4Mux_h
    port map (
            O => \N__27524\,
            I => \N__27515\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__27521\,
            I => \N__27512\
        );

    \I__4329\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27509\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__27515\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__4327\ : Odrv4
    port map (
            O => \N__27512\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__27509\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__4325\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27499\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__27499\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__27496\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27493\,
            I => \N__27487\
        );

    \I__4321\ : InMux
    port map (
            O => \N__27492\,
            I => \N__27487\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__27487\,
            I => \N__27482\
        );

    \I__4319\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27477\
        );

    \I__4318\ : InMux
    port map (
            O => \N__27485\,
            I => \N__27477\
        );

    \I__4317\ : Span4Mux_h
    port map (
            O => \N__27482\,
            I => \N__27474\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__27477\,
            I => \N__27471\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__27474\,
            I => \N__27468\
        );

    \I__4314\ : Span12Mux_v
    port map (
            O => \N__27471\,
            I => \N__27465\
        );

    \I__4313\ : Odrv4
    port map (
            O => \N__27468\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__4312\ : Odrv12
    port map (
            O => \N__27465\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__27460\,
            I => \N__27457\
        );

    \I__4310\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27454\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__27454\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__27451\,
            I => \N__27448\
        );

    \I__4307\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27445\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N__27442\
        );

    \I__4305\ : Span4Mux_h
    port map (
            O => \N__27442\,
            I => \N__27439\
        );

    \I__4304\ : Odrv4
    port map (
            O => \N__27439\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__27436\,
            I => \N__27433\
        );

    \I__4302\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27429\
        );

    \I__4301\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27426\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__27429\,
            I => \N__27423\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__27426\,
            I => \N__27419\
        );

    \I__4298\ : Span4Mux_v
    port map (
            O => \N__27423\,
            I => \N__27415\
        );

    \I__4297\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27412\
        );

    \I__4296\ : Span4Mux_v
    port map (
            O => \N__27419\,
            I => \N__27409\
        );

    \I__4295\ : InMux
    port map (
            O => \N__27418\,
            I => \N__27406\
        );

    \I__4294\ : Span4Mux_h
    port map (
            O => \N__27415\,
            I => \N__27401\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__27412\,
            I => \N__27401\
        );

    \I__4292\ : Odrv4
    port map (
            O => \N__27409\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__27406\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4290\ : Odrv4
    port map (
            O => \N__27401\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4289\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27391\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__27391\,
            I => \N__27388\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__27388\,
            I => \current_shift_inst.PI_CTRL.integrator_i_23\
        );

    \I__4286\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27382\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__27382\,
            I => \N__27379\
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__27379\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__27376\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__4282\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27370\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__27370\,
            I => \N__27367\
        );

    \I__4280\ : Odrv4
    port map (
            O => \N__27367\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__4279\ : InMux
    port map (
            O => \N__27364\,
            I => \N__27361\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__27361\,
            I => \N__27358\
        );

    \I__4277\ : Span4Mux_h
    port map (
            O => \N__27358\,
            I => \N__27355\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__27355\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__27352\,
            I => \N__27349\
        );

    \I__4274\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27345\
        );

    \I__4273\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27342\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__27345\,
            I => \N__27339\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__27342\,
            I => \N__27336\
        );

    \I__4270\ : Span4Mux_v
    port map (
            O => \N__27339\,
            I => \N__27331\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__27336\,
            I => \N__27328\
        );

    \I__4268\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27325\
        );

    \I__4267\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27322\
        );

    \I__4266\ : Span4Mux_v
    port map (
            O => \N__27331\,
            I => \N__27319\
        );

    \I__4265\ : Span4Mux_h
    port map (
            O => \N__27328\,
            I => \N__27314\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__27325\,
            I => \N__27314\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__27322\,
            I => \N__27311\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__27319\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__27314\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__4260\ : Odrv12
    port map (
            O => \N__27311\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__4259\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27300\
        );

    \I__4258\ : InMux
    port map (
            O => \N__27303\,
            I => \N__27296\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__27300\,
            I => \N__27293\
        );

    \I__4256\ : InMux
    port map (
            O => \N__27299\,
            I => \N__27290\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__27296\,
            I => \N__27287\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__27293\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__27290\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__4252\ : Odrv12
    port map (
            O => \N__27287\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__4251\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27276\
        );

    \I__4250\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27273\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__27276\,
            I => \N__27268\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__27273\,
            I => \N__27268\
        );

    \I__4247\ : Span4Mux_v
    port map (
            O => \N__27268\,
            I => \N__27263\
        );

    \I__4246\ : InMux
    port map (
            O => \N__27267\,
            I => \N__27260\
        );

    \I__4245\ : InMux
    port map (
            O => \N__27266\,
            I => \N__27257\
        );

    \I__4244\ : Span4Mux_h
    port map (
            O => \N__27263\,
            I => \N__27252\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__27260\,
            I => \N__27252\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__27257\,
            I => \N__27249\
        );

    \I__4241\ : Span4Mux_v
    port map (
            O => \N__27252\,
            I => \N__27246\
        );

    \I__4240\ : Span4Mux_v
    port map (
            O => \N__27249\,
            I => \N__27243\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__27246\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__4238\ : Odrv4
    port map (
            O => \N__27243\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__4237\ : CascadeMux
    port map (
            O => \N__27238\,
            I => \N__27235\
        );

    \I__4236\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27229\
        );

    \I__4235\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27229\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__27229\,
            I => \N__27226\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__27226\,
            I => \N__27222\
        );

    \I__4232\ : InMux
    port map (
            O => \N__27225\,
            I => \N__27219\
        );

    \I__4231\ : Odrv4
    port map (
            O => \N__27222\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__27219\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__4229\ : InMux
    port map (
            O => \N__27214\,
            I => \N__27211\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__27211\,
            I => \N__27208\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__27208\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__4226\ : InMux
    port map (
            O => \N__27205\,
            I => \bfn_11_10_0_\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__27202\,
            I => \N__27199\
        );

    \I__4224\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27196\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__27196\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__4222\ : CascadeMux
    port map (
            O => \N__27193\,
            I => \N__27190\
        );

    \I__4221\ : InMux
    port map (
            O => \N__27190\,
            I => \N__27186\
        );

    \I__4220\ : InMux
    port map (
            O => \N__27189\,
            I => \N__27182\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__27186\,
            I => \N__27179\
        );

    \I__4218\ : InMux
    port map (
            O => \N__27185\,
            I => \N__27176\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__27182\,
            I => \N__27172\
        );

    \I__4216\ : Span4Mux_v
    port map (
            O => \N__27179\,
            I => \N__27167\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__27176\,
            I => \N__27167\
        );

    \I__4214\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27164\
        );

    \I__4213\ : Odrv4
    port map (
            O => \N__27172\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__27167\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__27164\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__27157\,
            I => \N__27154\
        );

    \I__4209\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27151\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__27151\,
            I => \current_shift_inst.PI_CTRL.integrator_i_29\
        );

    \I__4207\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27144\
        );

    \I__4206\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27141\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__27144\,
            I => \N__27137\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__27141\,
            I => \N__27134\
        );

    \I__4203\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27130\
        );

    \I__4202\ : Span4Mux_v
    port map (
            O => \N__27137\,
            I => \N__27125\
        );

    \I__4201\ : Span4Mux_v
    port map (
            O => \N__27134\,
            I => \N__27125\
        );

    \I__4200\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27122\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__27130\,
            I => \N__27119\
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__27125\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__27122\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__27119\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__27112\,
            I => \N__27109\
        );

    \I__4194\ : InMux
    port map (
            O => \N__27109\,
            I => \N__27106\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__27106\,
            I => \current_shift_inst.PI_CTRL.integrator_i_28\
        );

    \I__4192\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27100\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__27100\,
            I => \N__27097\
        );

    \I__4190\ : Odrv12
    port map (
            O => \N__27097\,
            I => \current_shift_inst.PI_CTRL.integrator_i_11\
        );

    \I__4189\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27089\
        );

    \I__4188\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27084\
        );

    \I__4187\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27084\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__27089\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__27084\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\
        );

    \I__4184\ : InMux
    port map (
            O => \N__27079\,
            I => \N__27076\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__27076\,
            I => \current_shift_inst.PI_CTRL.integrator_i_25\
        );

    \I__4182\ : InMux
    port map (
            O => \N__27073\,
            I => \N__27070\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__27070\,
            I => \N__27067\
        );

    \I__4180\ : Odrv4
    port map (
            O => \N__27067\,
            I => \current_shift_inst.PI_CTRL.integrator_i_26\
        );

    \I__4179\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27061\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__27061\,
            I => \N__27058\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__27058\,
            I => \N__27055\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__27055\,
            I => \N__27052\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__27052\,
            I => \il_min_comp1_D1\
        );

    \I__4174\ : InMux
    port map (
            O => \N__27049\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\
        );

    \I__4173\ : InMux
    port map (
            O => \N__27046\,
            I => \N__27043\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__27043\,
            I => \N__27040\
        );

    \I__4171\ : Odrv4
    port map (
            O => \N__27040\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__4170\ : InMux
    port map (
            O => \N__27037\,
            I => \bfn_11_9_0_\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__27034\,
            I => \N__27031\
        );

    \I__4168\ : InMux
    port map (
            O => \N__27031\,
            I => \N__27028\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__27028\,
            I => \N__27025\
        );

    \I__4166\ : Odrv4
    port map (
            O => \N__27025\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__4165\ : InMux
    port map (
            O => \N__27022\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\
        );

    \I__4164\ : InMux
    port map (
            O => \N__27019\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\
        );

    \I__4163\ : InMux
    port map (
            O => \N__27016\,
            I => \N__27013\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__27013\,
            I => \N__27010\
        );

    \I__4161\ : Odrv4
    port map (
            O => \N__27010\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__4160\ : InMux
    port map (
            O => \N__27007\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__27004\,
            I => \N__27001\
        );

    \I__4158\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26998\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__26998\,
            I => \N__26995\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__26995\,
            I => \N__26992\
        );

    \I__4155\ : Odrv4
    port map (
            O => \N__26992\,
            I => \current_shift_inst.PI_CTRL.integrator_i_27\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26986\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__26986\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26983\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26980\,
            I => \N__26977\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__26977\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__4149\ : InMux
    port map (
            O => \N__26974\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\
        );

    \I__4148\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26968\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__26968\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26965\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__26962\,
            I => \N__26959\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26956\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__26956\,
            I => \N__26953\
        );

    \I__4142\ : Span4Mux_h
    port map (
            O => \N__26953\,
            I => \N__26950\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__26950\,
            I => \current_shift_inst.PI_CTRL.integrator_i_30\
        );

    \I__4140\ : CascadeMux
    port map (
            O => \N__26947\,
            I => \N__26944\
        );

    \I__4139\ : InMux
    port map (
            O => \N__26944\,
            I => \N__26941\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26941\,
            I => \N__26938\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__26938\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26935\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\
        );

    \I__4135\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26929\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26929\,
            I => \current_shift_inst.PI_CTRL.integrator_i_14\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__26926\,
            I => \N__26923\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26920\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__26920\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__4130\ : InMux
    port map (
            O => \N__26917\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26911\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__26911\,
            I => \N__26908\
        );

    \I__4127\ : Odrv4
    port map (
            O => \N__26908\,
            I => \current_shift_inst.PI_CTRL.integrator_i_15\
        );

    \I__4126\ : CascadeMux
    port map (
            O => \N__26905\,
            I => \N__26902\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26899\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__26899\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__4123\ : InMux
    port map (
            O => \N__26896\,
            I => \bfn_11_8_0_\
        );

    \I__4122\ : InMux
    port map (
            O => \N__26893\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\
        );

    \I__4121\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26887\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__26887\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__4119\ : InMux
    port map (
            O => \N__26884\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\
        );

    \I__4118\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26878\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__26878\,
            I => \N__26875\
        );

    \I__4116\ : Span4Mux_h
    port map (
            O => \N__26875\,
            I => \N__26872\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__26872\,
            I => \current_shift_inst.PI_CTRL.integrator_i_18\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__26869\,
            I => \N__26866\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26863\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__26863\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__4111\ : InMux
    port map (
            O => \N__26860\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__26857\,
            I => \N__26854\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26851\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__26851\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__4107\ : InMux
    port map (
            O => \N__26848\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\
        );

    \I__4106\ : InMux
    port map (
            O => \N__26845\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\
        );

    \I__4105\ : InMux
    port map (
            O => \N__26842\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__26839\,
            I => \N__26836\
        );

    \I__4103\ : InMux
    port map (
            O => \N__26836\,
            I => \N__26833\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26833\,
            I => \N__26830\
        );

    \I__4101\ : Odrv12
    port map (
            O => \N__26830\,
            I => \current_shift_inst.PI_CTRL.integrator_i_22\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__26827\,
            I => \N__26824\
        );

    \I__4099\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26821\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__26821\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26815\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__26815\,
            I => \N__26812\
        );

    \I__4095\ : Span4Mux_h
    port map (
            O => \N__26812\,
            I => \N__26809\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__26809\,
            I => \current_shift_inst.PI_CTRL.integrator_i_6\
        );

    \I__4093\ : InMux
    port map (
            O => \N__26806\,
            I => \N__26803\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__26803\,
            I => \N__26800\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__26800\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26797\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26791\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__26791\,
            I => \N__26788\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__26788\,
            I => \N__26785\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__26785\,
            I => \current_shift_inst.PI_CTRL.integrator_i_7\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26782\,
            I => \bfn_11_7_0_\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26779\,
            I => \N__26776\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__26776\,
            I => \N__26773\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__26773\,
            I => \current_shift_inst.PI_CTRL.integrator_i_8\
        );

    \I__4081\ : InMux
    port map (
            O => \N__26770\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\
        );

    \I__4080\ : InMux
    port map (
            O => \N__26767\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\
        );

    \I__4079\ : InMux
    port map (
            O => \N__26764\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\
        );

    \I__4078\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26758\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__26758\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__4076\ : InMux
    port map (
            O => \N__26755\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26749\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26746\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__26746\,
            I => \current_shift_inst.PI_CTRL.integrator_i_12\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__26743\,
            I => \N__26740\
        );

    \I__4071\ : InMux
    port map (
            O => \N__26740\,
            I => \N__26737\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__26737\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__4069\ : InMux
    port map (
            O => \N__26734\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\
        );

    \I__4068\ : InMux
    port map (
            O => \N__26731\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\
        );

    \I__4067\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26725\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__26725\,
            I => \N__26722\
        );

    \I__4065\ : Odrv12
    port map (
            O => \N__26722\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\
        );

    \I__4064\ : InMux
    port map (
            O => \N__26719\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\
        );

    \I__4063\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26713\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__26713\,
            I => \N__26710\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__26710\,
            I => \current_shift_inst.PI_CTRL.integrator_i_1\
        );

    \I__4060\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26704\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__26704\,
            I => \N__26701\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__26701\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\
        );

    \I__4057\ : InMux
    port map (
            O => \N__26698\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\
        );

    \I__4056\ : InMux
    port map (
            O => \N__26695\,
            I => \N__26692\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__26692\,
            I => \current_shift_inst.PI_CTRL.integrator_i_2\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26686\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26686\,
            I => \N__26683\
        );

    \I__4052\ : Odrv12
    port map (
            O => \N__26683\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__4051\ : InMux
    port map (
            O => \N__26680\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\
        );

    \I__4050\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26674\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__26674\,
            I => \N__26671\
        );

    \I__4048\ : Odrv4
    port map (
            O => \N__26671\,
            I => \current_shift_inst.PI_CTRL.integrator_i_3\
        );

    \I__4047\ : CascadeMux
    port map (
            O => \N__26668\,
            I => \N__26665\
        );

    \I__4046\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26662\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__26662\,
            I => \N__26659\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__26659\,
            I => \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7\
        );

    \I__4043\ : InMux
    port map (
            O => \N__26656\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\
        );

    \I__4042\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26650\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__26650\,
            I => \current_shift_inst.PI_CTRL.integrator_i_4\
        );

    \I__4040\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26644\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__26644\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__4038\ : InMux
    port map (
            O => \N__26641\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__26638\,
            I => \N__26635\
        );

    \I__4036\ : InMux
    port map (
            O => \N__26635\,
            I => \N__26632\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__26632\,
            I => \current_shift_inst.PI_CTRL.integrator_i_5\
        );

    \I__4034\ : CascadeMux
    port map (
            O => \N__26629\,
            I => \N__26626\
        );

    \I__4033\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26623\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__26623\,
            I => \N__26620\
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__26620\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__4030\ : InMux
    port map (
            O => \N__26617\,
            I => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\
        );

    \I__4029\ : InMux
    port map (
            O => \N__26614\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__4028\ : InMux
    port map (
            O => \N__26611\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__4027\ : InMux
    port map (
            O => \N__26608\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__4026\ : InMux
    port map (
            O => \N__26605\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__4025\ : InMux
    port map (
            O => \N__26602\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__4024\ : InMux
    port map (
            O => \N__26599\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__4023\ : InMux
    port map (
            O => \N__26596\,
            I => \bfn_10_24_0_\
        );

    \I__4022\ : InMux
    port map (
            O => \N__26593\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__4021\ : InMux
    port map (
            O => \N__26590\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__4020\ : InMux
    port map (
            O => \N__26587\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__4019\ : InMux
    port map (
            O => \N__26584\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__4018\ : InMux
    port map (
            O => \N__26581\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26578\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__4016\ : InMux
    port map (
            O => \N__26575\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__4015\ : InMux
    port map (
            O => \N__26572\,
            I => \bfn_10_25_0_\
        );

    \I__4014\ : InMux
    port map (
            O => \N__26569\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__4013\ : InMux
    port map (
            O => \N__26566\,
            I => \bfn_10_23_0_\
        );

    \I__4012\ : InMux
    port map (
            O => \N__26563\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__4011\ : InMux
    port map (
            O => \N__26560\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__4010\ : InMux
    port map (
            O => \N__26557\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26554\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26551\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__4007\ : InMux
    port map (
            O => \N__26548\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__4006\ : InMux
    port map (
            O => \N__26545\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26538\
        );

    \I__4004\ : CascadeMux
    port map (
            O => \N__26541\,
            I => \N__26535\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__26538\,
            I => \N__26532\
        );

    \I__4002\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26529\
        );

    \I__4001\ : Span4Mux_v
    port map (
            O => \N__26532\,
            I => \N__26526\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__26529\,
            I => \N__26523\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__26526\,
            I => \N__26520\
        );

    \I__3998\ : Span4Mux_v
    port map (
            O => \N__26523\,
            I => \N__26517\
        );

    \I__3997\ : Odrv4
    port map (
            O => \N__26520\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__26517\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__3995\ : InMux
    port map (
            O => \N__26512\,
            I => \N__26509\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__26509\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__3993\ : InMux
    port map (
            O => \N__26506\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__3992\ : InMux
    port map (
            O => \N__26503\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__3991\ : InMux
    port map (
            O => \N__26500\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__3990\ : InMux
    port map (
            O => \N__26497\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__3989\ : InMux
    port map (
            O => \N__26494\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__3988\ : InMux
    port map (
            O => \N__26491\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__26488\,
            I => \N__26485\
        );

    \I__3986\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26482\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__26482\,
            I => \N__26478\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__26481\,
            I => \N__26475\
        );

    \I__3983\ : Span4Mux_h
    port map (
            O => \N__26478\,
            I => \N__26470\
        );

    \I__3982\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26467\
        );

    \I__3981\ : InMux
    port map (
            O => \N__26474\,
            I => \N__26464\
        );

    \I__3980\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26461\
        );

    \I__3979\ : Span4Mux_h
    port map (
            O => \N__26470\,
            I => \N__26456\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__26467\,
            I => \N__26456\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__26464\,
            I => \N__26451\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__26461\,
            I => \N__26451\
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__26456\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__3974\ : Odrv12
    port map (
            O => \N__26451\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26443\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__26443\,
            I => \N__26439\
        );

    \I__3971\ : InMux
    port map (
            O => \N__26442\,
            I => \N__26435\
        );

    \I__3970\ : Span4Mux_h
    port map (
            O => \N__26439\,
            I => \N__26432\
        );

    \I__3969\ : InMux
    port map (
            O => \N__26438\,
            I => \N__26429\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__26435\,
            I => \N__26426\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__26432\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__26429\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__3965\ : Odrv4
    port map (
            O => \N__26426\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__3964\ : InMux
    port map (
            O => \N__26419\,
            I => \N__26416\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__26416\,
            I => \N__26412\
        );

    \I__3962\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26409\
        );

    \I__3961\ : Span4Mux_h
    port map (
            O => \N__26412\,
            I => \N__26406\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__26409\,
            I => \N__26403\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__26406\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__26403\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__26398\,
            I => \N__26395\
        );

    \I__3956\ : InMux
    port map (
            O => \N__26395\,
            I => \N__26392\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__26392\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__26389\,
            I => \N__26386\
        );

    \I__3953\ : InMux
    port map (
            O => \N__26386\,
            I => \N__26383\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__26383\,
            I => \N__26380\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__26380\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__3950\ : InMux
    port map (
            O => \N__26377\,
            I => \N__26373\
        );

    \I__3949\ : InMux
    port map (
            O => \N__26376\,
            I => \N__26370\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__26373\,
            I => \N__26365\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__26370\,
            I => \N__26362\
        );

    \I__3946\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26359\
        );

    \I__3945\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26356\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__26365\,
            I => \N__26349\
        );

    \I__3943\ : Span4Mux_v
    port map (
            O => \N__26362\,
            I => \N__26349\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__26359\,
            I => \N__26349\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__26356\,
            I => \N__26346\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__26349\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__3939\ : Odrv12
    port map (
            O => \N__26346\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__3938\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26338\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__26338\,
            I => \N__26334\
        );

    \I__3936\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26331\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__26334\,
            I => \N__26325\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__26331\,
            I => \N__26325\
        );

    \I__3933\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26322\
        );

    \I__3932\ : Span4Mux_v
    port map (
            O => \N__26325\,
            I => \N__26319\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__26322\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__26319\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__26314\,
            I => \N__26311\
        );

    \I__3928\ : InMux
    port map (
            O => \N__26311\,
            I => \N__26307\
        );

    \I__3927\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26304\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__26307\,
            I => \N__26299\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__26304\,
            I => \N__26296\
        );

    \I__3924\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26293\
        );

    \I__3923\ : InMux
    port map (
            O => \N__26302\,
            I => \N__26290\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__26299\,
            I => \N__26287\
        );

    \I__3921\ : Span4Mux_h
    port map (
            O => \N__26296\,
            I => \N__26282\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__26293\,
            I => \N__26282\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__26290\,
            I => \N__26279\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__26287\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__26282\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__3916\ : Odrv12
    port map (
            O => \N__26279\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__3915\ : CascadeMux
    port map (
            O => \N__26272\,
            I => \N__26269\
        );

    \I__3914\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26266\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__26266\,
            I => \N__26262\
        );

    \I__3912\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26259\
        );

    \I__3911\ : Span4Mux_v
    port map (
            O => \N__26262\,
            I => \N__26255\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__26259\,
            I => \N__26252\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26249\
        );

    \I__3908\ : Span4Mux_h
    port map (
            O => \N__26255\,
            I => \N__26244\
        );

    \I__3907\ : Span4Mux_v
    port map (
            O => \N__26252\,
            I => \N__26244\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__26249\,
            I => \N__26241\
        );

    \I__3905\ : Odrv4
    port map (
            O => \N__26244\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__3904\ : Odrv12
    port map (
            O => \N__26241\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__26236\,
            I => \N__26233\
        );

    \I__3902\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26230\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__26230\,
            I => \N__26227\
        );

    \I__3900\ : Odrv12
    port map (
            O => \N__26227\,
            I => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\
        );

    \I__3899\ : InMux
    port map (
            O => \N__26224\,
            I => \N__26220\
        );

    \I__3898\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26217\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__26220\,
            I => \N__26214\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__26217\,
            I => \N__26211\
        );

    \I__3895\ : Span4Mux_v
    port map (
            O => \N__26214\,
            I => \N__26208\
        );

    \I__3894\ : Span4Mux_v
    port map (
            O => \N__26211\,
            I => \N__26203\
        );

    \I__3893\ : Span4Mux_h
    port map (
            O => \N__26208\,
            I => \N__26200\
        );

    \I__3892\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26195\
        );

    \I__3891\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26195\
        );

    \I__3890\ : Span4Mux_h
    port map (
            O => \N__26203\,
            I => \N__26190\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__26200\,
            I => \N__26190\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__26195\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__3887\ : Odrv4
    port map (
            O => \N__26190\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__3886\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26182\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__26182\,
            I => \N__26177\
        );

    \I__3884\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26174\
        );

    \I__3883\ : InMux
    port map (
            O => \N__26180\,
            I => \N__26171\
        );

    \I__3882\ : Sp12to4
    port map (
            O => \N__26177\,
            I => \N__26164\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__26174\,
            I => \N__26164\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__26171\,
            I => \N__26164\
        );

    \I__3879\ : Span12Mux_v
    port map (
            O => \N__26164\,
            I => \N__26161\
        );

    \I__3878\ : Odrv12
    port map (
            O => \N__26161\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__3877\ : IoInMux
    port map (
            O => \N__26158\,
            I => \N__26155\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__26155\,
            I => \N__26152\
        );

    \I__3875\ : Span4Mux_s3_v
    port map (
            O => \N__26152\,
            I => \N__26149\
        );

    \I__3874\ : Span4Mux_h
    port map (
            O => \N__26149\,
            I => \N__26146\
        );

    \I__3873\ : Span4Mux_v
    port map (
            O => \N__26146\,
            I => \N__26143\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__26143\,
            I => \delay_measurement_inst.delay_hc_timer.N_397_i\
        );

    \I__3871\ : InMux
    port map (
            O => \N__26140\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__26137\,
            I => \N__26134\
        );

    \I__3869\ : InMux
    port map (
            O => \N__26134\,
            I => \N__26129\
        );

    \I__3868\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26126\
        );

    \I__3867\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26123\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__26129\,
            I => \N__26118\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__26126\,
            I => \N__26118\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__26123\,
            I => \N__26113\
        );

    \I__3863\ : Span4Mux_v
    port map (
            O => \N__26118\,
            I => \N__26113\
        );

    \I__3862\ : Span4Mux_v
    port map (
            O => \N__26113\,
            I => \N__26109\
        );

    \I__3861\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26106\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__26109\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__26106\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__3858\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26098\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__26098\,
            I => \N__26095\
        );

    \I__3856\ : Span4Mux_h
    port map (
            O => \N__26095\,
            I => \N__26090\
        );

    \I__3855\ : InMux
    port map (
            O => \N__26094\,
            I => \N__26087\
        );

    \I__3854\ : InMux
    port map (
            O => \N__26093\,
            I => \N__26084\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__26090\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__26087\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__26084\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__26077\,
            I => \N__26073\
        );

    \I__3849\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26070\
        );

    \I__3848\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26067\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26060\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__26067\,
            I => \N__26060\
        );

    \I__3845\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26057\
        );

    \I__3844\ : InMux
    port map (
            O => \N__26065\,
            I => \N__26054\
        );

    \I__3843\ : Span4Mux_v
    port map (
            O => \N__26060\,
            I => \N__26051\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__26057\,
            I => \N__26048\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__26054\,
            I => \N__26045\
        );

    \I__3840\ : Span4Mux_v
    port map (
            O => \N__26051\,
            I => \N__26042\
        );

    \I__3839\ : Span4Mux_h
    port map (
            O => \N__26048\,
            I => \N__26037\
        );

    \I__3838\ : Span4Mux_v
    port map (
            O => \N__26045\,
            I => \N__26037\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__26042\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__3836\ : Odrv4
    port map (
            O => \N__26037\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__3835\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__26029\,
            I => \N__26025\
        );

    \I__3833\ : InMux
    port map (
            O => \N__26028\,
            I => \N__26022\
        );

    \I__3832\ : Span4Mux_v
    port map (
            O => \N__26025\,
            I => \N__26018\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__26022\,
            I => \N__26015\
        );

    \I__3830\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26012\
        );

    \I__3829\ : Span4Mux_h
    port map (
            O => \N__26018\,
            I => \N__26009\
        );

    \I__3828\ : Span4Mux_v
    port map (
            O => \N__26015\,
            I => \N__26006\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__26012\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__26009\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__26006\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25996\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__25996\,
            I => \N__25991\
        );

    \I__3822\ : InMux
    port map (
            O => \N__25995\,
            I => \N__25988\
        );

    \I__3821\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25985\
        );

    \I__3820\ : Span4Mux_h
    port map (
            O => \N__25991\,
            I => \N__25980\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25988\,
            I => \N__25980\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__25985\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__25980\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__25975\,
            I => \N__25972\
        );

    \I__3815\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25968\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__25971\,
            I => \N__25965\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__25968\,
            I => \N__25962\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25959\
        );

    \I__3811\ : Span4Mux_v
    port map (
            O => \N__25962\,
            I => \N__25953\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__25959\,
            I => \N__25953\
        );

    \I__3809\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25949\
        );

    \I__3808\ : Span4Mux_h
    port map (
            O => \N__25953\,
            I => \N__25946\
        );

    \I__3807\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25943\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__25949\,
            I => \N__25940\
        );

    \I__3805\ : Span4Mux_v
    port map (
            O => \N__25946\,
            I => \N__25937\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__25943\,
            I => \N__25934\
        );

    \I__3803\ : Span4Mux_v
    port map (
            O => \N__25940\,
            I => \N__25931\
        );

    \I__3802\ : Odrv4
    port map (
            O => \N__25937\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__3801\ : Odrv4
    port map (
            O => \N__25934\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__25931\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25924\,
            I => \N__25919\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25923\,
            I => \N__25916\
        );

    \I__3797\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25912\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__25919\,
            I => \N__25909\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__25916\,
            I => \N__25906\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25915\,
            I => \N__25903\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__25912\,
            I => \N__25900\
        );

    \I__3792\ : Span4Mux_h
    port map (
            O => \N__25909\,
            I => \N__25897\
        );

    \I__3791\ : Span12Mux_v
    port map (
            O => \N__25906\,
            I => \N__25894\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__25903\,
            I => \N__25891\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__25900\,
            I => \N__25888\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__25897\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__3787\ : Odrv12
    port map (
            O => \N__25894\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__25891\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__3785\ : Odrv4
    port map (
            O => \N__25888\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__25879\,
            I => \N__25876\
        );

    \I__3783\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25872\
        );

    \I__3782\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25868\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__25872\,
            I => \N__25865\
        );

    \I__3780\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25862\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__25868\,
            I => \N__25859\
        );

    \I__3778\ : Span4Mux_h
    port map (
            O => \N__25865\,
            I => \N__25854\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__25862\,
            I => \N__25854\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__25859\,
            I => \N__25851\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__25854\,
            I => \N__25848\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__25851\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__3773\ : Odrv4
    port map (
            O => \N__25848\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__3772\ : InMux
    port map (
            O => \N__25843\,
            I => \N__25840\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__25840\,
            I => \N__25837\
        );

    \I__3770\ : Span4Mux_h
    port map (
            O => \N__25837\,
            I => \N__25834\
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__25834\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__3768\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25828\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__25828\,
            I => \N__25822\
        );

    \I__3766\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25819\
        );

    \I__3765\ : InMux
    port map (
            O => \N__25826\,
            I => \N__25816\
        );

    \I__3764\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25813\
        );

    \I__3763\ : Span4Mux_h
    port map (
            O => \N__25822\,
            I => \N__25808\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__25819\,
            I => \N__25808\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__25816\,
            I => \N__25803\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__25813\,
            I => \N__25803\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__25808\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__3758\ : Odrv12
    port map (
            O => \N__25803\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__3757\ : InMux
    port map (
            O => \N__25798\,
            I => \N__25795\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__25795\,
            I => \N__25791\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25787\
        );

    \I__3754\ : Span4Mux_h
    port map (
            O => \N__25791\,
            I => \N__25784\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25781\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__25787\,
            I => \N__25778\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__25784\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__25781\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__3749\ : Odrv12
    port map (
            O => \N__25778\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__25771\,
            I => \N__25768\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25768\,
            I => \N__25765\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__25765\,
            I => \N__25762\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__25762\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__3744\ : InMux
    port map (
            O => \N__25759\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25753\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__25753\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25750\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__25747\,
            I => \N__25744\
        );

    \I__3739\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25741\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__25741\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__3737\ : InMux
    port map (
            O => \N__25738\,
            I => \bfn_10_16_0_\
        );

    \I__3736\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25732\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__25732\,
            I => \N__25729\
        );

    \I__3734\ : Odrv12
    port map (
            O => \N__25729\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__3733\ : InMux
    port map (
            O => \N__25726\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__25723\,
            I => \N__25720\
        );

    \I__3731\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25717\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__25717\,
            I => \N__25714\
        );

    \I__3729\ : Odrv12
    port map (
            O => \N__25714\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__3728\ : InMux
    port map (
            O => \N__25711\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__3727\ : InMux
    port map (
            O => \N__25708\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__25705\,
            I => \N__25702\
        );

    \I__3725\ : InMux
    port map (
            O => \N__25702\,
            I => \N__25699\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__25699\,
            I => \N__25696\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__25696\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__3722\ : InMux
    port map (
            O => \N__25693\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__3721\ : InMux
    port map (
            O => \N__25690\,
            I => \N__25687\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25687\,
            I => \N__25684\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__25684\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__3718\ : InMux
    port map (
            O => \N__25681\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__25678\,
            I => \N__25675\
        );

    \I__3716\ : InMux
    port map (
            O => \N__25675\,
            I => \N__25672\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__25672\,
            I => \N__25669\
        );

    \I__3714\ : Span4Mux_h
    port map (
            O => \N__25669\,
            I => \N__25666\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__25666\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__3712\ : InMux
    port map (
            O => \N__25663\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__25660\,
            I => \N__25657\
        );

    \I__3710\ : InMux
    port map (
            O => \N__25657\,
            I => \N__25654\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__25654\,
            I => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25651\,
            I => \N__25648\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__25648\,
            I => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__25645\,
            I => \N__25642\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25639\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__25639\,
            I => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\
        );

    \I__3703\ : InMux
    port map (
            O => \N__25636\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__3702\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25630\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__25630\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__3700\ : InMux
    port map (
            O => \N__25627\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__3699\ : InMux
    port map (
            O => \N__25624\,
            I => \N__25621\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__25621\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__25618\,
            I => \N__25615\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25612\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__25612\,
            I => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\
        );

    \I__3694\ : InMux
    port map (
            O => \N__25609\,
            I => \N__25606\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__25606\,
            I => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__25603\,
            I => \N__25600\
        );

    \I__3691\ : InMux
    port map (
            O => \N__25600\,
            I => \N__25597\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__25597\,
            I => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\
        );

    \I__3689\ : InMux
    port map (
            O => \N__25594\,
            I => \N__25591\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__25591\,
            I => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\
        );

    \I__3687\ : CascadeMux
    port map (
            O => \N__25588\,
            I => \N__25585\
        );

    \I__3686\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25582\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__25582\,
            I => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\
        );

    \I__3684\ : InMux
    port map (
            O => \N__25579\,
            I => \N__25576\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__25576\,
            I => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\
        );

    \I__3682\ : CascadeMux
    port map (
            O => \N__25573\,
            I => \N__25570\
        );

    \I__3681\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25567\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__25567\,
            I => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\
        );

    \I__3679\ : InMux
    port map (
            O => \N__25564\,
            I => \N__25561\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__25561\,
            I => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__25558\,
            I => \N__25547\
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__25557\,
            I => \N__25543\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__25556\,
            I => \N__25539\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__25555\,
            I => \N__25535\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__25554\,
            I => \N__25532\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__25553\,
            I => \N__25528\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__25552\,
            I => \N__25524\
        );

    \I__3670\ : CascadeMux
    port map (
            O => \N__25551\,
            I => \N__25520\
        );

    \I__3669\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25501\
        );

    \I__3668\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25501\
        );

    \I__3667\ : InMux
    port map (
            O => \N__25546\,
            I => \N__25501\
        );

    \I__3666\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25501\
        );

    \I__3665\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25501\
        );

    \I__3664\ : InMux
    port map (
            O => \N__25539\,
            I => \N__25501\
        );

    \I__3663\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25501\
        );

    \I__3662\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25501\
        );

    \I__3661\ : InMux
    port map (
            O => \N__25532\,
            I => \N__25484\
        );

    \I__3660\ : InMux
    port map (
            O => \N__25531\,
            I => \N__25484\
        );

    \I__3659\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25484\
        );

    \I__3658\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25484\
        );

    \I__3657\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25484\
        );

    \I__3656\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25484\
        );

    \I__3655\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25484\
        );

    \I__3654\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25484\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__25518\,
            I => \N__25481\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__25501\,
            I => \N__25475\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__25484\,
            I => \N__25475\
        );

    \I__3650\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25470\
        );

    \I__3649\ : InMux
    port map (
            O => \N__25480\,
            I => \N__25470\
        );

    \I__3648\ : Span4Mux_v
    port map (
            O => \N__25475\,
            I => \N__25467\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__25470\,
            I => \N__25464\
        );

    \I__3646\ : Odrv4
    port map (
            O => \N__25467\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__3645\ : Odrv12
    port map (
            O => \N__25464\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25456\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__25456\,
            I => \N__25453\
        );

    \I__3642\ : Span4Mux_h
    port map (
            O => \N__25453\,
            I => \N__25450\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__25450\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__25447\,
            I => \N__25444\
        );

    \I__3639\ : InMux
    port map (
            O => \N__25444\,
            I => \N__25441\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__25441\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25438\,
            I => \N__25435\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__25435\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__25432\,
            I => \N__25429\
        );

    \I__3634\ : InMux
    port map (
            O => \N__25429\,
            I => \N__25426\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__25426\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__25423\,
            I => \N__25420\
        );

    \I__3631\ : InMux
    port map (
            O => \N__25420\,
            I => \N__25417\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__25417\,
            I => \N__25414\
        );

    \I__3629\ : Odrv12
    port map (
            O => \N__25414\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__3628\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25408\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__25408\,
            I => \N__25405\
        );

    \I__3626\ : Odrv4
    port map (
            O => \N__25405\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__3625\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25399\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__25399\,
            I => \N__25396\
        );

    \I__3623\ : Odrv12
    port map (
            O => \N__25396\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__3622\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25390\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__25390\,
            I => \N__25387\
        );

    \I__3620\ : Odrv12
    port map (
            O => \N__25387\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3619\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25381\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__25381\,
            I => \N__25376\
        );

    \I__3617\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25372\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__25379\,
            I => \N__25369\
        );

    \I__3615\ : Span4Mux_h
    port map (
            O => \N__25376\,
            I => \N__25366\
        );

    \I__3614\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25363\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__25372\,
            I => \N__25360\
        );

    \I__3612\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25357\
        );

    \I__3611\ : Span4Mux_v
    port map (
            O => \N__25366\,
            I => \N__25350\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__25363\,
            I => \N__25350\
        );

    \I__3609\ : Span4Mux_v
    port map (
            O => \N__25360\,
            I => \N__25350\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__25357\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__25350\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__3606\ : InMux
    port map (
            O => \N__25345\,
            I => \N__25333\
        );

    \I__3605\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25333\
        );

    \I__3604\ : InMux
    port map (
            O => \N__25343\,
            I => \N__25333\
        );

    \I__3603\ : InMux
    port map (
            O => \N__25342\,
            I => \N__25333\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__25333\,
            I => \N__25304\
        );

    \I__3601\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25295\
        );

    \I__3600\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25295\
        );

    \I__3599\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25295\
        );

    \I__3598\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25295\
        );

    \I__3597\ : InMux
    port map (
            O => \N__25328\,
            I => \N__25286\
        );

    \I__3596\ : InMux
    port map (
            O => \N__25327\,
            I => \N__25286\
        );

    \I__3595\ : InMux
    port map (
            O => \N__25326\,
            I => \N__25286\
        );

    \I__3594\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25286\
        );

    \I__3593\ : InMux
    port map (
            O => \N__25324\,
            I => \N__25277\
        );

    \I__3592\ : InMux
    port map (
            O => \N__25323\,
            I => \N__25277\
        );

    \I__3591\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25277\
        );

    \I__3590\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25277\
        );

    \I__3589\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25272\
        );

    \I__3588\ : InMux
    port map (
            O => \N__25319\,
            I => \N__25272\
        );

    \I__3587\ : InMux
    port map (
            O => \N__25318\,
            I => \N__25263\
        );

    \I__3586\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25263\
        );

    \I__3585\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25263\
        );

    \I__3584\ : InMux
    port map (
            O => \N__25315\,
            I => \N__25263\
        );

    \I__3583\ : InMux
    port map (
            O => \N__25314\,
            I => \N__25254\
        );

    \I__3582\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25254\
        );

    \I__3581\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25254\
        );

    \I__3580\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25254\
        );

    \I__3579\ : InMux
    port map (
            O => \N__25310\,
            I => \N__25245\
        );

    \I__3578\ : InMux
    port map (
            O => \N__25309\,
            I => \N__25245\
        );

    \I__3577\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25245\
        );

    \I__3576\ : InMux
    port map (
            O => \N__25307\,
            I => \N__25245\
        );

    \I__3575\ : Span4Mux_h
    port map (
            O => \N__25304\,
            I => \N__25240\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__25295\,
            I => \N__25240\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25235\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__25277\,
            I => \N__25235\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__25272\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__25263\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__25254\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__25245\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__25240\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__25235\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__3565\ : IoInMux
    port map (
            O => \N__25222\,
            I => \N__25219\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__25219\,
            I => \N__25216\
        );

    \I__3563\ : Span4Mux_s2_v
    port map (
            O => \N__25216\,
            I => \N__25213\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__25213\,
            I => s4_phy_c
        );

    \I__3561\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25207\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__25207\,
            I => \il_max_comp1_D1\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__25204\,
            I => \N__25201\
        );

    \I__3558\ : InMux
    port map (
            O => \N__25201\,
            I => \N__25198\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__25198\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__3556\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25192\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__25192\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__25189\,
            I => \N__25186\
        );

    \I__3553\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25183\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__25183\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__3551\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25177\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25174\
        );

    \I__3549\ : Odrv4
    port map (
            O => \N__25174\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__25171\,
            I => \N__25168\
        );

    \I__3547\ : InMux
    port map (
            O => \N__25168\,
            I => \N__25165\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__25165\,
            I => \N__25162\
        );

    \I__3545\ : Span4Mux_v
    port map (
            O => \N__25162\,
            I => \N__25159\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__25159\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__3543\ : InMux
    port map (
            O => \N__25156\,
            I => \N__25153\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__25153\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__25150\,
            I => \N__25147\
        );

    \I__3540\ : InMux
    port map (
            O => \N__25147\,
            I => \N__25144\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__25144\,
            I => \N__25141\
        );

    \I__3538\ : Span4Mux_v
    port map (
            O => \N__25141\,
            I => \N__25138\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__25138\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__3536\ : InMux
    port map (
            O => \N__25135\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__3535\ : IoInMux
    port map (
            O => \N__25132\,
            I => \N__25129\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__25129\,
            I => \N__25126\
        );

    \I__3533\ : Span12Mux_s3_v
    port map (
            O => \N__25126\,
            I => \N__25123\
        );

    \I__3532\ : Odrv12
    port map (
            O => \N__25123\,
            I => s3_phy_c
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__25120\,
            I => \N__25117\
        );

    \I__3530\ : InMux
    port map (
            O => \N__25117\,
            I => \N__25114\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__25114\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__3528\ : InMux
    port map (
            O => \N__25111\,
            I => \N__25108\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__25108\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__25105\,
            I => \N__25102\
        );

    \I__3525\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25099\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__25099\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__3523\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25093\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__25093\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__3521\ : InMux
    port map (
            O => \N__25090\,
            I => \N__25087\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__25087\,
            I => \N__25084\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__25084\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__25081\,
            I => \N__25078\
        );

    \I__3517\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25075\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__25075\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__3515\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25069\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__25069\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__25066\,
            I => \N__25063\
        );

    \I__3512\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25060\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__25060\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__3510\ : InMux
    port map (
            O => \N__25057\,
            I => \N__25054\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__25054\,
            I => \N__25051\
        );

    \I__3508\ : Odrv4
    port map (
            O => \N__25051\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__25048\,
            I => \N__25045\
        );

    \I__3506\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25042\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__25042\,
            I => \N__25039\
        );

    \I__3504\ : Odrv4
    port map (
            O => \N__25039\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__25036\,
            I => \N__25033\
        );

    \I__3502\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25030\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__25027\
        );

    \I__3500\ : Odrv12
    port map (
            O => \N__25027\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__3499\ : InMux
    port map (
            O => \N__25024\,
            I => \N__25021\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__25021\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__3497\ : InMux
    port map (
            O => \N__25018\,
            I => \N__25015\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__25015\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__25012\,
            I => \N__25009\
        );

    \I__3494\ : InMux
    port map (
            O => \N__25009\,
            I => \N__25006\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__25003\
        );

    \I__3492\ : Odrv4
    port map (
            O => \N__25003\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__3491\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24997\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__24997\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__24994\,
            I => \N__24991\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24991\,
            I => \N__24988\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__24988\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24982\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__24982\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__24979\,
            I => \N__24976\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24973\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__24973\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__3481\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24967\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__24967\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__24964\,
            I => \N__24961\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24958\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__24958\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__3476\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24946\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24954\,
            I => \N__24946\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24946\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__3472\ : Span4Mux_v
    port map (
            O => \N__24943\,
            I => \N__24939\
        );

    \I__3471\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24936\
        );

    \I__3470\ : Span4Mux_v
    port map (
            O => \N__24939\,
            I => \N__24933\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__24936\,
            I => \N__24930\
        );

    \I__3468\ : Odrv4
    port map (
            O => \N__24933\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__3467\ : Odrv12
    port map (
            O => \N__24930\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__24925\,
            I => \N__24922\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24916\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24916\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24916\,
            I => \N__24912\
        );

    \I__3462\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24909\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__24912\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24909\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__24904\,
            I => \N__24901\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24896\
        );

    \I__3457\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24891\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24899\,
            I => \N__24891\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__24896\,
            I => \N__24888\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__24891\,
            I => \N__24885\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__24888\,
            I => \N__24881\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__24885\,
            I => \N__24878\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24884\,
            I => \N__24875\
        );

    \I__3450\ : Span4Mux_v
    port map (
            O => \N__24881\,
            I => \N__24872\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__24878\,
            I => \N__24869\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__24875\,
            I => \N__24866\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__24872\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__24869\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__3445\ : Odrv12
    port map (
            O => \N__24866\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__24859\,
            I => \N__24855\
        );

    \I__3443\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24851\
        );

    \I__3442\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24848\
        );

    \I__3441\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24845\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__24851\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__24848\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__24845\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__24838\,
            I => \N__24835\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24830\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24834\,
            I => \N__24827\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24824\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__24830\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__24827\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__24824\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24817\,
            I => \N__24814\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__24814\,
            I => \N__24809\
        );

    \I__3428\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24806\
        );

    \I__3427\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24803\
        );

    \I__3426\ : Span4Mux_v
    port map (
            O => \N__24809\,
            I => \N__24795\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__24806\,
            I => \N__24795\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24803\,
            I => \N__24795\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24792\
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__24795\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__24792\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24783\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__24786\,
            I => \N__24779\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__24783\,
            I => \N__24776\
        );

    \I__3417\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24771\
        );

    \I__3416\ : InMux
    port map (
            O => \N__24779\,
            I => \N__24771\
        );

    \I__3415\ : Span4Mux_v
    port map (
            O => \N__24776\,
            I => \N__24768\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24771\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__24768\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24757\
        );

    \I__3411\ : InMux
    port map (
            O => \N__24762\,
            I => \N__24757\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__24757\,
            I => \N__24753\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24756\,
            I => \N__24749\
        );

    \I__3408\ : Sp12to4
    port map (
            O => \N__24753\,
            I => \N__24746\
        );

    \I__3407\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24743\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__24749\,
            I => \N__24740\
        );

    \I__3405\ : Span12Mux_v
    port map (
            O => \N__24746\,
            I => \N__24737\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__24743\,
            I => \N__24734\
        );

    \I__3403\ : Span4Mux_v
    port map (
            O => \N__24740\,
            I => \N__24731\
        );

    \I__3402\ : Odrv12
    port map (
            O => \N__24737\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__24734\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__24731\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__24724\,
            I => \N__24720\
        );

    \I__3398\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24715\
        );

    \I__3397\ : InMux
    port map (
            O => \N__24720\,
            I => \N__24715\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__24715\,
            I => \N__24712\
        );

    \I__3395\ : Span4Mux_h
    port map (
            O => \N__24712\,
            I => \N__24708\
        );

    \I__3394\ : InMux
    port map (
            O => \N__24711\,
            I => \N__24705\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__24708\,
            I => \N__24701\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__24705\,
            I => \N__24698\
        );

    \I__3391\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24695\
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__24701\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__24698\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__24695\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__24688\,
            I => \N__24684\
        );

    \I__3386\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24680\
        );

    \I__3385\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24675\
        );

    \I__3384\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24675\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__24680\,
            I => \N__24672\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__24675\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__3381\ : Odrv12
    port map (
            O => \N__24672\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24664\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__24664\,
            I => \N__24661\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__24661\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__3377\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24655\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__24655\,
            I => \N__24652\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__24652\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__3374\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24646\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24643\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__24643\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__3371\ : InMux
    port map (
            O => \N__24640\,
            I => \N__24637\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__24637\,
            I => \N__24634\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__24634\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__3368\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24628\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__24628\,
            I => \N__24625\
        );

    \I__3366\ : Span4Mux_v
    port map (
            O => \N__24625\,
            I => \N__24622\
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__24622\,
            I => \il_min_comp2_D1\
        );

    \I__3364\ : InMux
    port map (
            O => \N__24619\,
            I => \N__24616\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__24616\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\
        );

    \I__3362\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24610\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__24610\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__3360\ : InMux
    port map (
            O => \N__24607\,
            I => \N__24604\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__24604\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__3358\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24598\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__24598\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__3356\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24592\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__24592\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__3354\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24586\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__24586\,
            I => \N__24583\
        );

    \I__3352\ : Span12Mux_h
    port map (
            O => \N__24583\,
            I => \N__24580\
        );

    \I__3351\ : Odrv12
    port map (
            O => \N__24580\,
            I => il_max_comp1_c
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__24577\,
            I => \N__24574\
        );

    \I__3349\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24571\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__24571\,
            I => \N__24566\
        );

    \I__3347\ : InMux
    port map (
            O => \N__24570\,
            I => \N__24563\
        );

    \I__3346\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24560\
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__24566\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__24563\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__24560\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3342\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24550\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__24550\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__3340\ : InMux
    port map (
            O => \N__24547\,
            I => \N__24544\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__24544\,
            I => \current_shift_inst.PI_CTRL.un1_enablelt3_0\
        );

    \I__3338\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24538\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__24538\,
            I => \current_shift_inst.PI_CTRL.N_71\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__24535\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__24532\,
            I => \N__24529\
        );

    \I__3334\ : InMux
    port map (
            O => \N__24529\,
            I => \N__24526\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__24526\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__24523\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10_cascade_\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__24520\,
            I => \N__24517\
        );

    \I__3330\ : InMux
    port map (
            O => \N__24517\,
            I => \N__24514\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__24514\,
            I => \N__24511\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__24511\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__24508\,
            I => \N__24505\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24505\,
            I => \N__24500\
        );

    \I__3325\ : InMux
    port map (
            O => \N__24504\,
            I => \N__24497\
        );

    \I__3324\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24494\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__24500\,
            I => \N__24489\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__24497\,
            I => \N__24489\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__24494\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__24489\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__3319\ : InMux
    port map (
            O => \N__24484\,
            I => \bfn_8_24_0_\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__24481\,
            I => \N__24477\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__24480\,
            I => \N__24474\
        );

    \I__3316\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24470\
        );

    \I__3315\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24467\
        );

    \I__3314\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24464\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__24470\,
            I => \N__24459\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__24467\,
            I => \N__24459\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__24464\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__24459\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__3309\ : InMux
    port map (
            O => \N__24454\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__3308\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24444\
        );

    \I__3307\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24444\
        );

    \I__3306\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24441\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__24444\,
            I => \N__24438\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__24441\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__24438\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__3302\ : InMux
    port map (
            O => \N__24433\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__24430\,
            I => \N__24427\
        );

    \I__3300\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24422\
        );

    \I__3299\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24419\
        );

    \I__3298\ : InMux
    port map (
            O => \N__24425\,
            I => \N__24416\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24422\,
            I => \N__24411\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__24419\,
            I => \N__24411\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__24416\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__24411\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__3293\ : InMux
    port map (
            O => \N__24406\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__24403\,
            I => \N__24400\
        );

    \I__3291\ : InMux
    port map (
            O => \N__24400\,
            I => \N__24396\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24399\,
            I => \N__24393\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24396\,
            I => \N__24390\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__24393\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__24390\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__3286\ : InMux
    port map (
            O => \N__24385\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__3285\ : InMux
    port map (
            O => \N__24382\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__3284\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24376\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__24376\,
            I => \N__24372\
        );

    \I__3282\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24369\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__24372\,
            I => \N__24366\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__24369\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__24366\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__3278\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24358\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__24358\,
            I => \N__24355\
        );

    \I__3276\ : Odrv12
    port map (
            O => \N__24355\,
            I => il_min_comp1_c
        );

    \I__3275\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24345\
        );

    \I__3274\ : InMux
    port map (
            O => \N__24351\,
            I => \N__24345\
        );

    \I__3273\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24342\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__24345\,
            I => \N__24339\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__24342\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__24339\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__3269\ : InMux
    port map (
            O => \N__24334\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__24331\,
            I => \N__24328\
        );

    \I__3267\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24323\
        );

    \I__3266\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24320\
        );

    \I__3265\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24317\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__24323\,
            I => \N__24312\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__24320\,
            I => \N__24312\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__24317\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__24312\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__3260\ : InMux
    port map (
            O => \N__24307\,
            I => \bfn_8_23_0_\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__24304\,
            I => \N__24300\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__24303\,
            I => \N__24297\
        );

    \I__3257\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24293\
        );

    \I__3256\ : InMux
    port map (
            O => \N__24297\,
            I => \N__24290\
        );

    \I__3255\ : InMux
    port map (
            O => \N__24296\,
            I => \N__24287\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__24293\,
            I => \N__24282\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__24290\,
            I => \N__24282\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24287\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__24282\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__3250\ : InMux
    port map (
            O => \N__24277\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__3249\ : InMux
    port map (
            O => \N__24274\,
            I => \N__24267\
        );

    \I__3248\ : InMux
    port map (
            O => \N__24273\,
            I => \N__24267\
        );

    \I__3247\ : InMux
    port map (
            O => \N__24272\,
            I => \N__24264\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__24267\,
            I => \N__24261\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__24264\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__24261\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__3243\ : InMux
    port map (
            O => \N__24256\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__24253\,
            I => \N__24250\
        );

    \I__3241\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24245\
        );

    \I__3240\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24242\
        );

    \I__3239\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24239\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__24245\,
            I => \N__24234\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__24242\,
            I => \N__24234\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__24239\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__24234\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__3234\ : InMux
    port map (
            O => \N__24229\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__24226\,
            I => \N__24222\
        );

    \I__3232\ : InMux
    port map (
            O => \N__24225\,
            I => \N__24218\
        );

    \I__3231\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24215\
        );

    \I__3230\ : InMux
    port map (
            O => \N__24221\,
            I => \N__24212\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__24218\,
            I => \N__24207\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__24215\,
            I => \N__24207\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__24212\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__24207\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__3225\ : InMux
    port map (
            O => \N__24202\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__24199\,
            I => \N__24196\
        );

    \I__3223\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24191\
        );

    \I__3222\ : InMux
    port map (
            O => \N__24195\,
            I => \N__24188\
        );

    \I__3221\ : InMux
    port map (
            O => \N__24194\,
            I => \N__24185\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__24191\,
            I => \N__24180\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__24188\,
            I => \N__24180\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__24185\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__24180\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__3216\ : InMux
    port map (
            O => \N__24175\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__24172\,
            I => \N__24168\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__24171\,
            I => \N__24165\
        );

    \I__3213\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24159\
        );

    \I__3212\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24159\
        );

    \I__3211\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24156\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__24159\,
            I => \N__24153\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__24156\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__24153\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__3207\ : InMux
    port map (
            O => \N__24148\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__3206\ : InMux
    port map (
            O => \N__24145\,
            I => \N__24138\
        );

    \I__3205\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24138\
        );

    \I__3204\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24135\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__24138\,
            I => \N__24132\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__24135\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__24132\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__3200\ : InMux
    port map (
            O => \N__24127\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__3199\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24117\
        );

    \I__3198\ : InMux
    port map (
            O => \N__24123\,
            I => \N__24117\
        );

    \I__3197\ : InMux
    port map (
            O => \N__24122\,
            I => \N__24114\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__24117\,
            I => \N__24111\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__24114\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__24111\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__3193\ : InMux
    port map (
            O => \N__24106\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__24103\,
            I => \N__24100\
        );

    \I__3191\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24095\
        );

    \I__3190\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24092\
        );

    \I__3189\ : InMux
    port map (
            O => \N__24098\,
            I => \N__24089\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__24095\,
            I => \N__24084\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__24092\,
            I => \N__24084\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__24089\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__24084\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__3184\ : InMux
    port map (
            O => \N__24079\,
            I => \bfn_8_22_0_\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__24076\,
            I => \N__24072\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__24075\,
            I => \N__24069\
        );

    \I__3181\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24066\
        );

    \I__3180\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24062\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__24066\,
            I => \N__24059\
        );

    \I__3178\ : InMux
    port map (
            O => \N__24065\,
            I => \N__24056\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__24062\,
            I => \N__24051\
        );

    \I__3176\ : Span4Mux_h
    port map (
            O => \N__24059\,
            I => \N__24051\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__24056\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__24051\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__3173\ : InMux
    port map (
            O => \N__24046\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__3172\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24036\
        );

    \I__3171\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24036\
        );

    \I__3170\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24033\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__24036\,
            I => \N__24030\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__24033\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__24030\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__3166\ : InMux
    port map (
            O => \N__24025\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__24022\,
            I => \N__24019\
        );

    \I__3164\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24014\
        );

    \I__3163\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24011\
        );

    \I__3162\ : InMux
    port map (
            O => \N__24017\,
            I => \N__24008\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__24014\,
            I => \N__24003\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24003\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__24008\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__24003\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__3157\ : InMux
    port map (
            O => \N__23998\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__23995\,
            I => \N__23991\
        );

    \I__3155\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23987\
        );

    \I__3154\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23984\
        );

    \I__3153\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23981\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__23987\,
            I => \N__23976\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__23984\,
            I => \N__23976\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__23981\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__3149\ : Odrv4
    port map (
            O => \N__23976\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__3148\ : InMux
    port map (
            O => \N__23971\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__23968\,
            I => \N__23965\
        );

    \I__3146\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23960\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23957\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23954\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__23960\,
            I => \N__23949\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__23957\,
            I => \N__23949\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__23954\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__23949\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__3139\ : InMux
    port map (
            O => \N__23944\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__23941\,
            I => \N__23937\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__23940\,
            I => \N__23934\
        );

    \I__3136\ : InMux
    port map (
            O => \N__23937\,
            I => \N__23928\
        );

    \I__3135\ : InMux
    port map (
            O => \N__23934\,
            I => \N__23928\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23933\,
            I => \N__23925\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__23928\,
            I => \N__23922\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__23925\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__3131\ : Odrv4
    port map (
            O => \N__23922\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__3130\ : InMux
    port map (
            O => \N__23917\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23914\,
            I => \N__23909\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23906\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23903\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__23909\,
            I => \N__23900\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__23906\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__23903\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__23900\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23893\,
            I => \bfn_8_21_0_\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23887\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__23887\,
            I => \N__23882\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23879\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23876\
        );

    \I__3117\ : Span4Mux_v
    port map (
            O => \N__23882\,
            I => \N__23871\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23871\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__23876\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__3114\ : Odrv4
    port map (
            O => \N__23871\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23866\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__23863\,
            I => \N__23859\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__23862\,
            I => \N__23856\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23850\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23850\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23855\,
            I => \N__23847\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23850\,
            I => \N__23844\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__23847\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__23844\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__3104\ : InMux
    port map (
            O => \N__23839\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__23836\,
            I => \N__23832\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__23835\,
            I => \N__23829\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23823\
        );

    \I__3100\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23823\
        );

    \I__3099\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23820\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23823\,
            I => \N__23817\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__23820\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__23817\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__3095\ : InMux
    port map (
            O => \N__23812\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__23809\,
            I => \N__23806\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23801\
        );

    \I__3092\ : InMux
    port map (
            O => \N__23805\,
            I => \N__23798\
        );

    \I__3091\ : InMux
    port map (
            O => \N__23804\,
            I => \N__23795\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23801\,
            I => \N__23790\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23790\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__23795\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__23790\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23785\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__23782\,
            I => \N__23779\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23774\
        );

    \I__3083\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23771\
        );

    \I__3082\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23768\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__23774\,
            I => \N__23763\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__23771\,
            I => \N__23763\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__23768\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__3078\ : Odrv4
    port map (
            O => \N__23763\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__3077\ : InMux
    port map (
            O => \N__23758\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__23755\,
            I => \N__23752\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23748\
        );

    \I__3074\ : InMux
    port map (
            O => \N__23751\,
            I => \N__23745\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__23748\,
            I => \N__23739\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__23745\,
            I => \N__23739\
        );

    \I__3071\ : InMux
    port map (
            O => \N__23744\,
            I => \N__23736\
        );

    \I__3070\ : Span4Mux_h
    port map (
            O => \N__23739\,
            I => \N__23733\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__23736\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__23733\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__3067\ : InMux
    port map (
            O => \N__23728\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__3066\ : InMux
    port map (
            O => \N__23725\,
            I => \N__23722\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__23722\,
            I => \N__23719\
        );

    \I__3064\ : Span4Mux_v
    port map (
            O => \N__23719\,
            I => \N__23716\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__23716\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__3062\ : InMux
    port map (
            O => \N__23713\,
            I => \N__23710\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__23710\,
            I => \N__23707\
        );

    \I__3060\ : Span4Mux_v
    port map (
            O => \N__23707\,
            I => \N__23704\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__23704\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__23701\,
            I => \N__23698\
        );

    \I__3057\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23695\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__23695\,
            I => \N__23692\
        );

    \I__3055\ : Span4Mux_v
    port map (
            O => \N__23692\,
            I => \N__23689\
        );

    \I__3054\ : Odrv4
    port map (
            O => \N__23689\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__3053\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23683\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__23683\,
            I => \N__23680\
        );

    \I__3051\ : Odrv12
    port map (
            O => \N__23680\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__3050\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23674\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__23674\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__3048\ : InMux
    port map (
            O => \N__23671\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__3047\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23665\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__23665\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__3045\ : InMux
    port map (
            O => \N__23662\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__3044\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23656\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__23656\,
            I => \N__23653\
        );

    \I__3042\ : Odrv4
    port map (
            O => \N__23653\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23650\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__3040\ : InMux
    port map (
            O => \N__23647\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__23644\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\
        );

    \I__3038\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23638\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__23638\,
            I => \N__23635\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__23635\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__3035\ : InMux
    port map (
            O => \N__23632\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__3034\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23626\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__23626\,
            I => \N__23623\
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__23623\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__3031\ : InMux
    port map (
            O => \N__23620\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__3030\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23614\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__23614\,
            I => \N__23611\
        );

    \I__3028\ : Odrv4
    port map (
            O => \N__23611\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__3027\ : InMux
    port map (
            O => \N__23608\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__3026\ : InMux
    port map (
            O => \N__23605\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__3025\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23599\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__23599\,
            I => \N__23596\
        );

    \I__3023\ : Odrv4
    port map (
            O => \N__23596\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__3022\ : InMux
    port map (
            O => \N__23593\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23587\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__23587\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__3019\ : InMux
    port map (
            O => \N__23584\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__3018\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23578\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__23578\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__3016\ : InMux
    port map (
            O => \N__23575\,
            I => \bfn_8_16_0_\
        );

    \I__3015\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23569\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__23569\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__3013\ : InMux
    port map (
            O => \N__23566\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__3012\ : InMux
    port map (
            O => \N__23563\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__3011\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23557\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__23557\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23554\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__3008\ : InMux
    port map (
            O => \N__23551\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__3007\ : InMux
    port map (
            O => \N__23548\,
            I => \N__23545\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__23545\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23542\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__3004\ : InMux
    port map (
            O => \N__23539\,
            I => \N__23536\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__23536\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__3002\ : InMux
    port map (
            O => \N__23533\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23530\,
            I => \N__23527\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__23527\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__2999\ : InMux
    port map (
            O => \N__23524\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__2998\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23518\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__23518\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__2996\ : InMux
    port map (
            O => \N__23515\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__2995\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23509\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__23509\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__2993\ : InMux
    port map (
            O => \N__23506\,
            I => \bfn_8_15_0_\
        );

    \I__2992\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23500\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__23500\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__2990\ : InMux
    port map (
            O => \N__23497\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__2989\ : InMux
    port map (
            O => \N__23494\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__2988\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23488\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__23488\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__2986\ : InMux
    port map (
            O => \N__23485\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__2985\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23479\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__23479\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__2983\ : InMux
    port map (
            O => \N__23476\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__2982\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23470\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__23470\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__2980\ : InMux
    port map (
            O => \N__23467\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__2979\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23461\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__23461\,
            I => \N__23458\
        );

    \I__2977\ : Span4Mux_v
    port map (
            O => \N__23458\,
            I => \N__23455\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__23455\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__2975\ : InMux
    port map (
            O => \N__23452\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__2974\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23446\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__23446\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__2972\ : InMux
    port map (
            O => \N__23443\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__2971\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23437\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__23437\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__2969\ : InMux
    port map (
            O => \N__23434\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__2968\ : InMux
    port map (
            O => \N__23431\,
            I => \bfn_8_14_0_\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__23428\,
            I => \current_shift_inst.PI_CTRL.N_72_cascade_\
        );

    \I__2966\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23422\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__23422\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__2964\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23416\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__23416\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2962\ : InMux
    port map (
            O => \N__23413\,
            I => \N__23410\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__23410\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2960\ : InMux
    port map (
            O => \N__23407\,
            I => \N__23404\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__23404\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2958\ : InMux
    port map (
            O => \N__23401\,
            I => \N__23398\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__23398\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2956\ : InMux
    port map (
            O => \N__23395\,
            I => \N__23392\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__23392\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__23389\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__2953\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23383\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__23383\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__2951\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23377\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__23377\,
            I => \N__23374\
        );

    \I__2949\ : Span12Mux_h
    port map (
            O => \N__23374\,
            I => \N__23371\
        );

    \I__2948\ : Odrv12
    port map (
            O => \N__23371\,
            I => il_min_comp2_c
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__23368\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\
        );

    \I__2946\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23362\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__23362\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\
        );

    \I__2944\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23356\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__23356\,
            I => \N__23353\
        );

    \I__2942\ : Span4Mux_h
    port map (
            O => \N__23353\,
            I => \N__23350\
        );

    \I__2941\ : Odrv4
    port map (
            O => \N__23350\,
            I => \il_max_comp2_D1\
        );

    \I__2940\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23344\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__23344\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23338\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__23338\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__23335\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__23332\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__2934\ : InMux
    port map (
            O => \N__23329\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23326\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__2932\ : InMux
    port map (
            O => \N__23323\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__2931\ : InMux
    port map (
            O => \N__23320\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__2930\ : InMux
    port map (
            O => \N__23317\,
            I => \bfn_7_22_0_\
        );

    \I__2929\ : InMux
    port map (
            O => \N__23314\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__2928\ : InMux
    port map (
            O => \N__23311\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__2927\ : InMux
    port map (
            O => \N__23308\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__2926\ : InMux
    port map (
            O => \N__23305\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__2925\ : InMux
    port map (
            O => \N__23302\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__2924\ : InMux
    port map (
            O => \N__23299\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__2923\ : InMux
    port map (
            O => \N__23296\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__2922\ : InMux
    port map (
            O => \N__23293\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__2921\ : InMux
    port map (
            O => \N__23290\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__2920\ : InMux
    port map (
            O => \N__23287\,
            I => \bfn_7_21_0_\
        );

    \I__2919\ : InMux
    port map (
            O => \N__23284\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__2918\ : InMux
    port map (
            O => \N__23281\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__2917\ : InMux
    port map (
            O => \N__23278\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__2916\ : InMux
    port map (
            O => \N__23275\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__2915\ : InMux
    port map (
            O => \N__23272\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__2914\ : InMux
    port map (
            O => \N__23269\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__2913\ : InMux
    port map (
            O => \N__23266\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__2912\ : InMux
    port map (
            O => \N__23263\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__2911\ : InMux
    port map (
            O => \N__23260\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__2910\ : InMux
    port map (
            O => \N__23257\,
            I => \bfn_7_20_0_\
        );

    \I__2909\ : InMux
    port map (
            O => \N__23254\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__2908\ : InMux
    port map (
            O => \N__23251\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__2907\ : InMux
    port map (
            O => \N__23248\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__2906\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23241\
        );

    \I__2905\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23238\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__23241\,
            I => \N__23235\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__23238\,
            I => \N__23232\
        );

    \I__2902\ : Span4Mux_h
    port map (
            O => \N__23235\,
            I => \N__23227\
        );

    \I__2901\ : Span4Mux_h
    port map (
            O => \N__23232\,
            I => \N__23227\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__23227\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2899\ : InMux
    port map (
            O => \N__23224\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__23221\,
            I => \N__23217\
        );

    \I__2897\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23214\
        );

    \I__2896\ : InMux
    port map (
            O => \N__23217\,
            I => \N__23211\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__23214\,
            I => \N__23206\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__23211\,
            I => \N__23206\
        );

    \I__2893\ : Span4Mux_h
    port map (
            O => \N__23206\,
            I => \N__23203\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__23203\,
            I => \N__23200\
        );

    \I__2891\ : Odrv4
    port map (
            O => \N__23200\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2890\ : InMux
    port map (
            O => \N__23197\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2889\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23188\
        );

    \I__2888\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23188\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__23188\,
            I => \N__23185\
        );

    \I__2886\ : Odrv4
    port map (
            O => \N__23185\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2885\ : InMux
    port map (
            O => \N__23182\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2884\ : InMux
    port map (
            O => \N__23179\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2883\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23172\
        );

    \I__2882\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23162\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__23172\,
            I => \N__23159\
        );

    \I__2880\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23150\
        );

    \I__2879\ : InMux
    port map (
            O => \N__23170\,
            I => \N__23150\
        );

    \I__2878\ : InMux
    port map (
            O => \N__23169\,
            I => \N__23150\
        );

    \I__2877\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23150\
        );

    \I__2876\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23143\
        );

    \I__2875\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23143\
        );

    \I__2874\ : InMux
    port map (
            O => \N__23165\,
            I => \N__23143\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__23162\,
            I => \N__23139\
        );

    \I__2872\ : Span4Mux_s3_h
    port map (
            O => \N__23159\,
            I => \N__23136\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__23150\,
            I => \N__23133\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__23143\,
            I => \N__23130\
        );

    \I__2869\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23127\
        );

    \I__2868\ : Span4Mux_s3_h
    port map (
            O => \N__23139\,
            I => \N__23124\
        );

    \I__2867\ : Span4Mux_v
    port map (
            O => \N__23136\,
            I => \N__23119\
        );

    \I__2866\ : Span4Mux_s3_h
    port map (
            O => \N__23133\,
            I => \N__23119\
        );

    \I__2865\ : Span4Mux_h
    port map (
            O => \N__23130\,
            I => \N__23114\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__23127\,
            I => \N__23114\
        );

    \I__2863\ : Span4Mux_h
    port map (
            O => \N__23124\,
            I => \N__23111\
        );

    \I__2862\ : Span4Mux_h
    port map (
            O => \N__23119\,
            I => \N__23108\
        );

    \I__2861\ : Span4Mux_h
    port map (
            O => \N__23114\,
            I => \N__23105\
        );

    \I__2860\ : Odrv4
    port map (
            O => \N__23111\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__23108\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__23105\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2857\ : InMux
    port map (
            O => \N__23098\,
            I => \N__23095\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__23095\,
            I => \N__23091\
        );

    \I__2855\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23088\
        );

    \I__2854\ : Span4Mux_v
    port map (
            O => \N__23091\,
            I => \N__23085\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__23088\,
            I => \N__23082\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__23085\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2851\ : Odrv12
    port map (
            O => \N__23082\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2850\ : InMux
    port map (
            O => \N__23077\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__2848\ : InMux
    port map (
            O => \N__23071\,
            I => \N__23067\
        );

    \I__2847\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23064\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__23067\,
            I => \N__23059\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__23064\,
            I => \N__23059\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__23059\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2843\ : InMux
    port map (
            O => \N__23056\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2842\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23049\
        );

    \I__2841\ : InMux
    port map (
            O => \N__23052\,
            I => \N__23046\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__23049\,
            I => \N__23043\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__23046\,
            I => \N__23040\
        );

    \I__2838\ : Span4Mux_h
    port map (
            O => \N__23043\,
            I => \N__23037\
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__23040\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__23037\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2835\ : InMux
    port map (
            O => \N__23032\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2834\ : InMux
    port map (
            O => \N__23029\,
            I => \N__23023\
        );

    \I__2833\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23023\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__23023\,
            I => \N__23020\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__23020\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2830\ : InMux
    port map (
            O => \N__23017\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2829\ : InMux
    port map (
            O => \N__23014\,
            I => \N__23008\
        );

    \I__2828\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23008\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__23008\,
            I => \N__23005\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__23005\,
            I => \N__23002\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__23002\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22999\,
            I => \bfn_7_12_0_\
        );

    \I__2823\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22990\
        );

    \I__2822\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22990\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__22987\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22984\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__22981\,
            I => \N__22977\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__22980\,
            I => \N__22974\
        );

    \I__2816\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22969\
        );

    \I__2815\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22969\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__22969\,
            I => \N__22966\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__22966\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22963\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__22960\,
            I => \N__22956\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22959\,
            I => \N__22951\
        );

    \I__2809\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22951\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__22948\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22945\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__22942\,
            I => \N__22938\
        );

    \I__2804\ : InMux
    port map (
            O => \N__22941\,
            I => \N__22935\
        );

    \I__2803\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22932\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__22935\,
            I => \N__22927\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__22932\,
            I => \N__22927\
        );

    \I__2800\ : Span4Mux_h
    port map (
            O => \N__22927\,
            I => \N__22924\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__22924\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2798\ : InMux
    port map (
            O => \N__22921\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22914\
        );

    \I__2796\ : InMux
    port map (
            O => \N__22917\,
            I => \N__22911\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__22914\,
            I => \N__22906\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__22911\,
            I => \N__22906\
        );

    \I__2793\ : Span4Mux_v
    port map (
            O => \N__22906\,
            I => \N__22903\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__22903\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2791\ : InMux
    port map (
            O => \N__22900\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__22897\,
            I => \N__22893\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__22896\,
            I => \N__22890\
        );

    \I__2788\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22885\
        );

    \I__2787\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22885\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__22885\,
            I => \N__22882\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__22882\,
            I => \N__22879\
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__22879\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2783\ : InMux
    port map (
            O => \N__22876\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2782\ : InMux
    port map (
            O => \N__22873\,
            I => \N__22867\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22867\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__22867\,
            I => \N__22864\
        );

    \I__2779\ : Span4Mux_h
    port map (
            O => \N__22864\,
            I => \N__22861\
        );

    \I__2778\ : Odrv4
    port map (
            O => \N__22861\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22858\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__22855\,
            I => \N__22852\
        );

    \I__2775\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22848\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22851\,
            I => \N__22845\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__22848\,
            I => \N__22842\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__22845\,
            I => \N__22839\
        );

    \I__2771\ : Span4Mux_v
    port map (
            O => \N__22842\,
            I => \N__22836\
        );

    \I__2770\ : Span4Mux_h
    port map (
            O => \N__22839\,
            I => \N__22833\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__22836\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__22833\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22828\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2766\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22821\
        );

    \I__2765\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22818\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__22821\,
            I => \N__22815\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__22818\,
            I => \N__22812\
        );

    \I__2762\ : Span4Mux_h
    port map (
            O => \N__22815\,
            I => \N__22809\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__22812\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__22809\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2759\ : InMux
    port map (
            O => \N__22804\,
            I => \bfn_7_11_0_\
        );

    \I__2758\ : InMux
    port map (
            O => \N__22801\,
            I => \N__22797\
        );

    \I__2757\ : InMux
    port map (
            O => \N__22800\,
            I => \N__22794\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__22797\,
            I => \N__22791\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__22794\,
            I => \N__22788\
        );

    \I__2754\ : Span4Mux_h
    port map (
            O => \N__22791\,
            I => \N__22785\
        );

    \I__2753\ : Odrv12
    port map (
            O => \N__22788\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2752\ : Odrv4
    port map (
            O => \N__22785\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2751\ : InMux
    port map (
            O => \N__22780\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22773\
        );

    \I__2749\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22770\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__22773\,
            I => \N__22767\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__22770\,
            I => \N__22764\
        );

    \I__2746\ : Span4Mux_h
    port map (
            O => \N__22767\,
            I => \N__22761\
        );

    \I__2745\ : Span4Mux_h
    port map (
            O => \N__22764\,
            I => \N__22758\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__22761\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__22758\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22753\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22750\,
            I => \N__22747\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__22747\,
            I => \N__22743\
        );

    \I__2739\ : InMux
    port map (
            O => \N__22746\,
            I => \N__22740\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__22743\,
            I => \N__22737\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__22740\,
            I => \N__22734\
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__22737\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__22734\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2734\ : InMux
    port map (
            O => \N__22729\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2733\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22721\
        );

    \I__2732\ : InMux
    port map (
            O => \N__22725\,
            I => \N__22716\
        );

    \I__2731\ : InMux
    port map (
            O => \N__22724\,
            I => \N__22716\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__22721\,
            I => \N__22713\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22710\
        );

    \I__2728\ : Span4Mux_h
    port map (
            O => \N__22713\,
            I => \N__22707\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__22710\,
            I => \N__22704\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__22707\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__22704\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2724\ : InMux
    port map (
            O => \N__22699\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2723\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22693\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__22693\,
            I => \N__22687\
        );

    \I__2721\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22684\
        );

    \I__2720\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22679\
        );

    \I__2719\ : InMux
    port map (
            O => \N__22690\,
            I => \N__22679\
        );

    \I__2718\ : Span4Mux_v
    port map (
            O => \N__22687\,
            I => \N__22676\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__22684\,
            I => \N__22671\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22671\
        );

    \I__2715\ : Span4Mux_h
    port map (
            O => \N__22676\,
            I => \N__22668\
        );

    \I__2714\ : Span4Mux_h
    port map (
            O => \N__22671\,
            I => \N__22665\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__22668\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__22665\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2711\ : InMux
    port map (
            O => \N__22660\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__2709\ : InMux
    port map (
            O => \N__22654\,
            I => \N__22651\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__22651\,
            I => \N__22647\
        );

    \I__2707\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22644\
        );

    \I__2706\ : Span4Mux_v
    port map (
            O => \N__22647\,
            I => \N__22641\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__22644\,
            I => \N__22637\
        );

    \I__2704\ : Span4Mux_s1_h
    port map (
            O => \N__22641\,
            I => \N__22634\
        );

    \I__2703\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22631\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__22637\,
            I => \N__22628\
        );

    \I__2701\ : Span4Mux_h
    port map (
            O => \N__22634\,
            I => \N__22623\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__22631\,
            I => \N__22623\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__22628\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__22623\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2697\ : InMux
    port map (
            O => \N__22618\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2696\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22612\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__22612\,
            I => \N__22609\
        );

    \I__2694\ : Span4Mux_s3_h
    port map (
            O => \N__22609\,
            I => \N__22604\
        );

    \I__2693\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22601\
        );

    \I__2692\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22598\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__22604\,
            I => \N__22593\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22593\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__22598\,
            I => \N__22590\
        );

    \I__2688\ : Span4Mux_h
    port map (
            O => \N__22593\,
            I => \N__22587\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__22590\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__22587\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2685\ : InMux
    port map (
            O => \N__22582\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__22579\,
            I => \N__22575\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__22578\,
            I => \N__22572\
        );

    \I__2682\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22568\
        );

    \I__2681\ : InMux
    port map (
            O => \N__22572\,
            I => \N__22565\
        );

    \I__2680\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22562\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__22568\,
            I => \N__22559\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__22565\,
            I => \N__22556\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__22562\,
            I => \N__22551\
        );

    \I__2676\ : Span4Mux_v
    port map (
            O => \N__22559\,
            I => \N__22551\
        );

    \I__2675\ : Odrv12
    port map (
            O => \N__22556\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2674\ : Odrv4
    port map (
            O => \N__22551\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2673\ : InMux
    port map (
            O => \N__22546\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2672\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22539\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__22542\,
            I => \N__22536\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__22539\,
            I => \N__22533\
        );

    \I__2669\ : InMux
    port map (
            O => \N__22536\,
            I => \N__22530\
        );

    \I__2668\ : Span4Mux_h
    port map (
            O => \N__22533\,
            I => \N__22525\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__22530\,
            I => \N__22525\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__22525\,
            I => \N__22521\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22524\,
            I => \N__22518\
        );

    \I__2664\ : Sp12to4
    port map (
            O => \N__22521\,
            I => \N__22513\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__22518\,
            I => \N__22513\
        );

    \I__2662\ : Odrv12
    port map (
            O => \N__22513\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2661\ : InMux
    port map (
            O => \N__22510\,
            I => \bfn_7_10_0_\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__22507\,
            I => \N__22504\
        );

    \I__2659\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22499\
        );

    \I__2658\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22496\
        );

    \I__2657\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22493\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22490\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__22496\,
            I => \N__22487\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__22493\,
            I => \N__22484\
        );

    \I__2653\ : Span4Mux_h
    port map (
            O => \N__22490\,
            I => \N__22479\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__22487\,
            I => \N__22479\
        );

    \I__2651\ : Odrv12
    port map (
            O => \N__22484\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__22479\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2649\ : InMux
    port map (
            O => \N__22474\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2648\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22465\
        );

    \I__2647\ : InMux
    port map (
            O => \N__22470\,
            I => \N__22465\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__22465\,
            I => \N__22462\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__22462\,
            I => \N__22459\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__22459\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2643\ : InMux
    port map (
            O => \N__22456\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2642\ : InMux
    port map (
            O => \N__22453\,
            I => \N__22450\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__22450\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2640\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22444\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__22444\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\
        );

    \I__2638\ : InMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__22438\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22432\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__2634\ : Span4Mux_s3_h
    port map (
            O => \N__22429\,
            I => \N__22426\
        );

    \I__2633\ : Span4Mux_h
    port map (
            O => \N__22426\,
            I => \N__22423\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__22423\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2631\ : InMux
    port map (
            O => \N__22420\,
            I => \N__22417\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__22417\,
            I => \N__22414\
        );

    \I__2629\ : Span12Mux_s7_h
    port map (
            O => \N__22414\,
            I => \N__22411\
        );

    \I__2628\ : Odrv12
    port map (
            O => \N__22411\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2627\ : InMux
    port map (
            O => \N__22408\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2626\ : InMux
    port map (
            O => \N__22405\,
            I => \N__22402\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__22402\,
            I => \N__22399\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__22399\,
            I => \N__22396\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__22396\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2622\ : InMux
    port map (
            O => \N__22393\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2621\ : InMux
    port map (
            O => \N__22390\,
            I => \N__22387\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__22387\,
            I => \N__22384\
        );

    \I__2619\ : Span4Mux_s1_h
    port map (
            O => \N__22384\,
            I => \N__22379\
        );

    \I__2618\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22376\
        );

    \I__2617\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22373\
        );

    \I__2616\ : Span4Mux_h
    port map (
            O => \N__22379\,
            I => \N__22370\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__22376\,
            I => pwm_duty_input_3
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__22373\,
            I => pwm_duty_input_3
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__22370\,
            I => pwm_duty_input_3
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__22363\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__22360\,
            I => \N__22352\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__22359\,
            I => \N__22349\
        );

    \I__2609\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22346\
        );

    \I__2608\ : InMux
    port map (
            O => \N__22357\,
            I => \N__22335\
        );

    \I__2607\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22335\
        );

    \I__2606\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22335\
        );

    \I__2605\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22335\
        );

    \I__2604\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22335\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__22346\,
            I => \N__22330\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__22335\,
            I => \N__22330\
        );

    \I__2601\ : Span4Mux_v
    port map (
            O => \N__22330\,
            I => \N__22326\
        );

    \I__2600\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22323\
        );

    \I__2599\ : Span4Mux_h
    port map (
            O => \N__22326\,
            I => \N__22320\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N__22317\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__22320\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__22317\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2595\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22309\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__22309\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2593\ : InMux
    port map (
            O => \N__22306\,
            I => \N__22303\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__22303\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2591\ : InMux
    port map (
            O => \N__22300\,
            I => \N__22297\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__22297\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22291\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__22291\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__2587\ : InMux
    port map (
            O => \N__22288\,
            I => \N__22285\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__22285\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2585\ : InMux
    port map (
            O => \N__22282\,
            I => \N__22279\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__22279\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2583\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22273\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__22273\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__22270\,
            I => \current_shift_inst.PI_CTRL.N_53_cascade_\
        );

    \I__2580\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22261\
        );

    \I__2579\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22261\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22258\
        );

    \I__2577\ : Span4Mux_h
    port map (
            O => \N__22258\,
            I => \N__22254\
        );

    \I__2576\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22251\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__22254\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__22251\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__2573\ : InMux
    port map (
            O => \N__22246\,
            I => \N__22243\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__22243\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__22240\,
            I => \N__22237\
        );

    \I__2570\ : InMux
    port map (
            O => \N__22237\,
            I => \N__22234\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__22234\,
            I => \current_shift_inst.PI_CTRL.N_155\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__22231\,
            I => \N__22227\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__22230\,
            I => \N__22224\
        );

    \I__2566\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22218\
        );

    \I__2565\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22218\
        );

    \I__2564\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22215\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__22218\,
            I => \N__22210\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__22215\,
            I => \N__22210\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__22210\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2560\ : ClkMux
    port map (
            O => \N__22207\,
            I => \N__22204\
        );

    \I__2559\ : GlobalMux
    port map (
            O => \N__22204\,
            I => \N__22201\
        );

    \I__2558\ : gio2CtrlBuf
    port map (
            O => \N__22201\,
            I => delay_hc_input_c_g
        );

    \I__2557\ : InMux
    port map (
            O => \N__22198\,
            I => \N__22195\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__22195\,
            I => \N__22192\
        );

    \I__2555\ : Odrv12
    port map (
            O => \N__22192\,
            I => il_max_comp2_c
        );

    \I__2554\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22186\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__22186\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__22183\,
            I => \N__22179\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__22182\,
            I => \N__22176\
        );

    \I__2550\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22169\
        );

    \I__2549\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22169\
        );

    \I__2548\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22166\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__22174\,
            I => \N__22163\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22160\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__22166\,
            I => \N__22157\
        );

    \I__2544\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22153\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__22160\,
            I => \N__22148\
        );

    \I__2542\ : Span4Mux_v
    port map (
            O => \N__22157\,
            I => \N__22148\
        );

    \I__2541\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22145\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__22153\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__22148\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__22145\,
            I => \current_shift_inst.PI_CTRL.N_153\
        );

    \I__2537\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22134\
        );

    \I__2536\ : InMux
    port map (
            O => \N__22137\,
            I => \N__22131\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__22134\,
            I => \N__22128\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__22131\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__22128\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__2532\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22115\
        );

    \I__2531\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22106\
        );

    \I__2530\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22106\
        );

    \I__2529\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22106\
        );

    \I__2528\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22106\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__22118\,
            I => \N__22103\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__22115\,
            I => \N__22100\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__22106\,
            I => \N__22097\
        );

    \I__2524\ : InMux
    port map (
            O => \N__22103\,
            I => \N__22092\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__22100\,
            I => \N__22089\
        );

    \I__2522\ : Span4Mux_h
    port map (
            O => \N__22097\,
            I => \N__22086\
        );

    \I__2521\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22081\
        );

    \I__2520\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22081\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__22092\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__22089\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__22086\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__22081\,
            I => \current_shift_inst.PI_CTRL.N_53\
        );

    \I__2515\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22069\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__22069\,
            I => \N__22066\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__22066\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__2512\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22060\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__22060\,
            I => \N__22055\
        );

    \I__2510\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22052\
        );

    \I__2509\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22049\
        );

    \I__2508\ : Span4Mux_h
    port map (
            O => \N__22055\,
            I => \N__22046\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__22052\,
            I => \N__22043\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__22049\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__22046\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__22043\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__22036\,
            I => \N__22033\
        );

    \I__2502\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22030\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__22030\,
            I => \N__22027\
        );

    \I__2500\ : Span4Mux_h
    port map (
            O => \N__22027\,
            I => \N__22023\
        );

    \I__2499\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22020\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__22023\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__22020\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__2496\ : CascadeMux
    port map (
            O => \N__22015\,
            I => \N__22010\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__22014\,
            I => \N__22006\
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__22013\,
            I => \N__22000\
        );

    \I__2493\ : InMux
    port map (
            O => \N__22010\,
            I => \N__21991\
        );

    \I__2492\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21991\
        );

    \I__2491\ : InMux
    port map (
            O => \N__22006\,
            I => \N__21991\
        );

    \I__2490\ : InMux
    port map (
            O => \N__22005\,
            I => \N__21988\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__22004\,
            I => \N__21985\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__22003\,
            I => \N__21982\
        );

    \I__2487\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21978\
        );

    \I__2486\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21975\
        );

    \I__2485\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21972\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__21991\,
            I => \N__21969\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__21988\,
            I => \N__21964\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21961\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21982\,
            I => \N__21958\
        );

    \I__2480\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21955\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21978\,
            I => \N__21948\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__21975\,
            I => \N__21948\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__21972\,
            I => \N__21948\
        );

    \I__2476\ : Span4Mux_v
    port map (
            O => \N__21969\,
            I => \N__21945\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21940\
        );

    \I__2474\ : InMux
    port map (
            O => \N__21967\,
            I => \N__21940\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__21964\,
            I => \N__21929\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__21961\,
            I => \N__21929\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21958\,
            I => \N__21929\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__21955\,
            I => \N__21929\
        );

    \I__2469\ : Span4Mux_h
    port map (
            O => \N__21948\,
            I => \N__21929\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__21945\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__21940\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__21929\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\
        );

    \I__2465\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21919\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__21919\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21916\,
            I => \N__21911\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21915\,
            I => \N__21908\
        );

    \I__2461\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21905\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__21911\,
            I => \N__21902\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__21908\,
            I => \N__21899\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21905\,
            I => \N__21896\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__21902\,
            I => \N__21893\
        );

    \I__2456\ : Span4Mux_h
    port map (
            O => \N__21899\,
            I => \N__21890\
        );

    \I__2455\ : Span4Mux_s1_h
    port map (
            O => \N__21896\,
            I => \N__21887\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__21893\,
            I => pwm_duty_input_9
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__21890\,
            I => pwm_duty_input_9
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__21887\,
            I => pwm_duty_input_9
        );

    \I__2451\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21875\
        );

    \I__2450\ : CascadeMux
    port map (
            O => \N__21879\,
            I => \N__21872\
        );

    \I__2449\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21869\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__21875\,
            I => \N__21866\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21863\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__21869\,
            I => \N__21860\
        );

    \I__2445\ : Span4Mux_h
    port map (
            O => \N__21866\,
            I => \N__21857\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__21863\,
            I => \N__21854\
        );

    \I__2443\ : Span4Mux_s2_h
    port map (
            O => \N__21860\,
            I => \N__21851\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__21857\,
            I => pwm_duty_input_6
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__21854\,
            I => pwm_duty_input_6
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__21851\,
            I => pwm_duty_input_6
        );

    \I__2439\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21841\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__21841\,
            I => \N__21836\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21840\,
            I => \N__21833\
        );

    \I__2436\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21830\
        );

    \I__2435\ : Span4Mux_v
    port map (
            O => \N__21836\,
            I => \N__21825\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__21833\,
            I => \N__21825\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__21830\,
            I => \N__21822\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__21825\,
            I => pwm_duty_input_8
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__21822\,
            I => pwm_duty_input_8
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__21817\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\
        );

    \I__2429\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21808\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21808\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__21808\,
            I => \N__21797\
        );

    \I__2426\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21794\
        );

    \I__2425\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21779\
        );

    \I__2424\ : InMux
    port map (
            O => \N__21805\,
            I => \N__21779\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21804\,
            I => \N__21779\
        );

    \I__2422\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21779\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21779\
        );

    \I__2420\ : InMux
    port map (
            O => \N__21801\,
            I => \N__21779\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21779\
        );

    \I__2418\ : Span4Mux_h
    port map (
            O => \N__21797\,
            I => \N__21774\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__21794\,
            I => \N__21774\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__21779\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__21774\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2414\ : InMux
    port map (
            O => \N__21769\,
            I => \N__21765\
        );

    \I__2413\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21762\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__21765\,
            I => \N__21756\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__21762\,
            I => \N__21756\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21753\
        );

    \I__2409\ : Span4Mux_s3_h
    port map (
            O => \N__21756\,
            I => \N__21750\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__21753\,
            I => \current_shift_inst.PI_CTRL.N_154\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__21750\,
            I => \current_shift_inst.PI_CTRL.N_154\
        );

    \I__2406\ : InMux
    port map (
            O => \N__21745\,
            I => \N__21741\
        );

    \I__2405\ : InMux
    port map (
            O => \N__21744\,
            I => \N__21738\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__21741\,
            I => \N__21735\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21730\
        );

    \I__2402\ : Span4Mux_v
    port map (
            O => \N__21735\,
            I => \N__21730\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__21730\,
            I => pwm_duty_input_2
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__21727\,
            I => \N__21724\
        );

    \I__2399\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21719\
        );

    \I__2398\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21716\
        );

    \I__2397\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21713\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21710\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21707\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__21713\,
            I => \N__21704\
        );

    \I__2393\ : Sp12to4
    port map (
            O => \N__21710\,
            I => \N__21699\
        );

    \I__2392\ : Span12Mux_v
    port map (
            O => \N__21707\,
            I => \N__21699\
        );

    \I__2391\ : Span4Mux_s1_h
    port map (
            O => \N__21704\,
            I => \N__21696\
        );

    \I__2390\ : Odrv12
    port map (
            O => \N__21699\,
            I => pwm_duty_input_7
        );

    \I__2389\ : Odrv4
    port map (
            O => \N__21696\,
            I => pwm_duty_input_7
        );

    \I__2388\ : InMux
    port map (
            O => \N__21691\,
            I => \N__21687\
        );

    \I__2387\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21683\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__21687\,
            I => \N__21680\
        );

    \I__2385\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21677\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__21683\,
            I => \N__21674\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__21680\,
            I => \N__21669\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__21677\,
            I => \N__21669\
        );

    \I__2381\ : Span4Mux_s1_h
    port map (
            O => \N__21674\,
            I => \N__21666\
        );

    \I__2380\ : Odrv4
    port map (
            O => \N__21669\,
            I => pwm_duty_input_5
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__21666\,
            I => pwm_duty_input_5
        );

    \I__2378\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21658\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__21658\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\
        );

    \I__2376\ : InMux
    port map (
            O => \N__21655\,
            I => \N__21652\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__21652\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__21649\,
            I => \N__21645\
        );

    \I__2373\ : InMux
    port map (
            O => \N__21648\,
            I => \N__21641\
        );

    \I__2372\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21638\
        );

    \I__2371\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21635\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__21641\,
            I => \N__21632\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__21638\,
            I => \N__21629\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__21635\,
            I => \N__21626\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__21632\,
            I => \N__21619\
        );

    \I__2366\ : Span4Mux_h
    port map (
            O => \N__21629\,
            I => \N__21619\
        );

    \I__2365\ : Span4Mux_v
    port map (
            O => \N__21626\,
            I => \N__21619\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__21619\,
            I => pwm_duty_input_4
        );

    \I__2363\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21613\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__21613\,
            I => \N__21610\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__21610\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__2360\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21583\
        );

    \I__2359\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21583\
        );

    \I__2358\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21583\
        );

    \I__2357\ : InMux
    port map (
            O => \N__21604\,
            I => \N__21583\
        );

    \I__2356\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21583\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21583\
        );

    \I__2354\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21583\
        );

    \I__2353\ : InMux
    port map (
            O => \N__21600\,
            I => \N__21580\
        );

    \I__2352\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21575\
        );

    \I__2351\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21575\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__21583\,
            I => \N__21568\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__21580\,
            I => \N__21568\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__21575\,
            I => \N__21568\
        );

    \I__2347\ : Span4Mux_v
    port map (
            O => \N__21568\,
            I => \N__21565\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__21565\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__21562\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__21559\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__21556\,
            I => \N__21553\
        );

    \I__2342\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21550\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__21550\,
            I => \N__21547\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__21547\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__21544\,
            I => \N__21541\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21538\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__21538\,
            I => \N__21535\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__21535\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__21532\,
            I => \N__21529\
        );

    \I__2334\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21526\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__21526\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__21523\,
            I => \N__21520\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21517\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__21517\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__2329\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21511\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__21511\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__2326\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21502\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__21502\,
            I => \N__21499\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__21499\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__2322\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21490\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__21490\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__21487\,
            I => \N__21484\
        );

    \I__2319\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21481\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__21481\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__2317\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21475\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__21475\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__21472\,
            I => \N__21469\
        );

    \I__2314\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21466\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__21466\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__21463\,
            I => \N__21460\
        );

    \I__2311\ : InMux
    port map (
            O => \N__21460\,
            I => \N__21457\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__21457\,
            I => \N__21454\
        );

    \I__2309\ : Span4Mux_h
    port map (
            O => \N__21454\,
            I => \N__21451\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__21451\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__21448\,
            I => \N__21445\
        );

    \I__2306\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21442\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__21442\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__2304\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21436\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__21436\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__21433\,
            I => \N__21425\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__21432\,
            I => \N__21420\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__21431\,
            I => \N__21415\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__21430\,
            I => \N__21412\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__21429\,
            I => \N__21403\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__21428\,
            I => \N__21400\
        );

    \I__2296\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21397\
        );

    \I__2295\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21382\
        );

    \I__2294\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21382\
        );

    \I__2293\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21382\
        );

    \I__2292\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21382\
        );

    \I__2291\ : InMux
    port map (
            O => \N__21418\,
            I => \N__21382\
        );

    \I__2290\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21382\
        );

    \I__2289\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21382\
        );

    \I__2288\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21379\
        );

    \I__2287\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21373\
        );

    \I__2286\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21373\
        );

    \I__2285\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21366\
        );

    \I__2284\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21366\
        );

    \I__2283\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21366\
        );

    \I__2282\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21361\
        );

    \I__2281\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21361\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__21397\,
            I => \N__21356\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__21382\,
            I => \N__21356\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__21379\,
            I => \N__21338\
        );

    \I__2277\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21335\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__21373\,
            I => \N__21330\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__21366\,
            I => \N__21330\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__21361\,
            I => \N__21325\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__21356\,
            I => \N__21325\
        );

    \I__2272\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21308\
        );

    \I__2271\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21308\
        );

    \I__2270\ : InMux
    port map (
            O => \N__21353\,
            I => \N__21308\
        );

    \I__2269\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21308\
        );

    \I__2268\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21308\
        );

    \I__2267\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21308\
        );

    \I__2266\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21308\
        );

    \I__2265\ : InMux
    port map (
            O => \N__21348\,
            I => \N__21308\
        );

    \I__2264\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21293\
        );

    \I__2263\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21293\
        );

    \I__2262\ : InMux
    port map (
            O => \N__21345\,
            I => \N__21293\
        );

    \I__2261\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21293\
        );

    \I__2260\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21293\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21293\
        );

    \I__2258\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21293\
        );

    \I__2257\ : Span12Mux_v
    port map (
            O => \N__21338\,
            I => \N__21286\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21286\
        );

    \I__2255\ : Span12Mux_s1_h
    port map (
            O => \N__21330\,
            I => \N__21286\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__21325\,
            I => \N_19_1\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__21308\,
            I => \N_19_1\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__21293\,
            I => \N_19_1\
        );

    \I__2251\ : Odrv12
    port map (
            O => \N__21286\,
            I => \N_19_1\
        );

    \I__2250\ : InMux
    port map (
            O => \N__21277\,
            I => \N__21274\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__21274\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__2248\ : InMux
    port map (
            O => \N__21271\,
            I => \N__21268\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__21268\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\
        );

    \I__2246\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21262\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__21262\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__2244\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21256\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__21256\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__2242\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21250\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__21250\,
            I => \N__21247\
        );

    \I__2240\ : Span4Mux_s2_h
    port map (
            O => \N__21247\,
            I => \N__21243\
        );

    \I__2239\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21240\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__21243\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__21240\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__21235\,
            I => \N__21232\
        );

    \I__2235\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21229\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__21229\,
            I => \N__21226\
        );

    \I__2233\ : Span4Mux_v
    port map (
            O => \N__21226\,
            I => \N__21223\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__21223\,
            I => \current_shift_inst.PI_CTRL.N_149\
        );

    \I__2231\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21217\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__21217\,
            I => \N__21213\
        );

    \I__2229\ : InMux
    port map (
            O => \N__21216\,
            I => \N__21210\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__21213\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__21210\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__2226\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21201\
        );

    \I__2225\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21198\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__21201\,
            I => \N__21192\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__21198\,
            I => \N__21192\
        );

    \I__2222\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21189\
        );

    \I__2221\ : Span4Mux_v
    port map (
            O => \N__21192\,
            I => \N__21186\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__21189\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__21186\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__2218\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21178\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__21178\,
            I => \N__21175\
        );

    \I__2216\ : Glb2LocalMux
    port map (
            O => \N__21175\,
            I => \N__21172\
        );

    \I__2215\ : GlobalMux
    port map (
            O => \N__21172\,
            I => clk_12mhz
        );

    \I__2214\ : IoInMux
    port map (
            O => \N__21169\,
            I => \N__21166\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__21166\,
            I => \N__21163\
        );

    \I__2212\ : Span4Mux_s0_v
    port map (
            O => \N__21163\,
            I => \N__21160\
        );

    \I__2211\ : Span4Mux_h
    port map (
            O => \N__21160\,
            I => \N__21157\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__21157\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2209\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21151\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__21151\,
            I => \N__21148\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__21148\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__21145\,
            I => \N__21142\
        );

    \I__2205\ : InMux
    port map (
            O => \N__21142\,
            I => \N__21139\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__21139\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__2203\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21133\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__21133\,
            I => \N__21130\
        );

    \I__2201\ : Span4Mux_h
    port map (
            O => \N__21130\,
            I => \N__21127\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__21127\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__2199\ : InMux
    port map (
            O => \N__21124\,
            I => \N__21121\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__21121\,
            I => \N__21118\
        );

    \I__2197\ : Odrv4
    port map (
            O => \N__21118\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1\
        );

    \I__2196\ : InMux
    port map (
            O => \N__21115\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__2195\ : InMux
    port map (
            O => \N__21112\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__2194\ : InMux
    port map (
            O => \N__21109\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__2193\ : InMux
    port map (
            O => \N__21106\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__2192\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21100\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__21100\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__2190\ : InMux
    port map (
            O => \N__21097\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__2189\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21091\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__21091\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__2187\ : InMux
    port map (
            O => \N__21088\,
            I => \bfn_3_10_0_\
        );

    \I__2186\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21082\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__21082\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__2184\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21076\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__21076\,
            I => \N__21073\
        );

    \I__2182\ : Span4Mux_h
    port map (
            O => \N__21073\,
            I => \N__21070\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__21070\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8\
        );

    \I__2180\ : InMux
    port map (
            O => \N__21067\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__2179\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21060\
        );

    \I__2178\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21057\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__21060\,
            I => \N__21054\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__21057\,
            I => \N__21051\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__21054\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__21051\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__21046\,
            I => \N__21042\
        );

    \I__2172\ : InMux
    port map (
            O => \N__21045\,
            I => \N__21038\
        );

    \I__2171\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21035\
        );

    \I__2170\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21032\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__21038\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__21035\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__21032\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2166\ : InMux
    port map (
            O => \N__21025\,
            I => \N__21022\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__21022\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__2164\ : InMux
    port map (
            O => \N__21019\,
            I => \N__21016\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__21016\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__2162\ : InMux
    port map (
            O => \N__21013\,
            I => \N__21008\
        );

    \I__2161\ : InMux
    port map (
            O => \N__21012\,
            I => \N__21005\
        );

    \I__2160\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21002\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__21008\,
            I => \N__20997\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__21005\,
            I => \N__20997\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__21002\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__20997\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20992\,
            I => \N__20989\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20989\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2153\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20981\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20978\
        );

    \I__2151\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20975\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__20981\,
            I => \N__20972\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__20978\,
            I => \N__20969\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__20975\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__20972\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__20969\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__20962\,
            I => \N__20959\
        );

    \I__2144\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20956\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__20956\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20953\,
            I => \N__20949\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20945\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20942\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20939\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__20945\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__20942\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__20939\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20929\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__20929\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2133\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20922\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20918\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__20922\,
            I => \N__20915\
        );

    \I__2130\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20912\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20918\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__20915\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__20912\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20905\,
            I => \N__20902\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20902\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2124\ : InMux
    port map (
            O => \N__20899\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2123\ : IoInMux
    port map (
            O => \N__20896\,
            I => \N__20893\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__20893\,
            I => \N__20890\
        );

    \I__2121\ : Span4Mux_s3_v
    port map (
            O => \N__20890\,
            I => \N__20887\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__20887\,
            I => \N__20884\
        );

    \I__2119\ : Sp12to4
    port map (
            O => \N__20884\,
            I => \N__20881\
        );

    \I__2118\ : Span12Mux_h
    port map (
            O => \N__20881\,
            I => \N__20878\
        );

    \I__2117\ : Odrv12
    port map (
            O => \N__20878\,
            I => pwm_output_c
        );

    \I__2116\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20872\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__20872\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20866\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__20866\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__2112\ : InMux
    port map (
            O => \N__20863\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__2111\ : InMux
    port map (
            O => \N__20860\,
            I => \N__20857\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__20857\,
            I => \N__20854\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__20854\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__2108\ : InMux
    port map (
            O => \N__20851\,
            I => \N__20848\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__20848\,
            I => \N__20845\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__20845\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20842\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20835\
        );

    \I__2103\ : InMux
    port map (
            O => \N__20838\,
            I => \N__20831\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__20835\,
            I => \N__20828\
        );

    \I__2101\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20825\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20831\,
            I => \N__20820\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__20828\,
            I => \N__20820\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__20825\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__20820\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20815\,
            I => \N__20812\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__20812\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2094\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20804\
        );

    \I__2093\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20801\
        );

    \I__2092\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20798\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__20804\,
            I => \N__20793\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__20801\,
            I => \N__20793\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__20798\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__20793\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20785\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__20785\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__20782\,
            I => \N__20779\
        );

    \I__2084\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20776\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__20776\,
            I => \N__20773\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__20773\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__2081\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20766\
        );

    \I__2080\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20763\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20766\,
            I => \N__20757\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__20763\,
            I => \N__20757\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20754\
        );

    \I__2076\ : Span4Mux_v
    port map (
            O => \N__20757\,
            I => \N__20751\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20754\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__20751\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2073\ : InMux
    port map (
            O => \N__20746\,
            I => \N__20743\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__20743\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20735\
        );

    \I__2070\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20732\
        );

    \I__2069\ : InMux
    port map (
            O => \N__20738\,
            I => \N__20729\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__20735\,
            I => \N__20724\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__20732\,
            I => \N__20724\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__20729\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__20724\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__20719\,
            I => \N__20716\
        );

    \I__2063\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__20713\,
            I => \N__20710\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__20710\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__2060\ : InMux
    port map (
            O => \N__20707\,
            I => \N__20704\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__20704\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2058\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20696\
        );

    \I__2057\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20693\
        );

    \I__2056\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20690\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__20696\,
            I => \N__20685\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__20693\,
            I => \N__20685\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__20690\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__20685\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2051\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20677\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__20677\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2049\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20669\
        );

    \I__2048\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20666\
        );

    \I__2047\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20663\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__20669\,
            I => \N__20658\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__20666\,
            I => \N__20658\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__20663\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__20658\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2042\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20650\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__20650\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2040\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__20644\,
            I => \N__20641\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__20641\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\
        );

    \I__2037\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20635\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__20635\,
            I => \N__20632\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__20632\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\
        );

    \I__2034\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20626\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__20626\,
            I => \N__20623\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__20623\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\
        );

    \I__2031\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20617\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__20617\,
            I => \N__20614\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__20614\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0\
        );

    \I__2028\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20608\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__20608\,
            I => \N__20605\
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__20605\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0\
        );

    \I__2025\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20599\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__20599\,
            I => \N__20596\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__20596\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0\
        );

    \I__2022\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20590\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__20590\,
            I => \N__20587\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__20587\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0\
        );

    \I__2019\ : InMux
    port map (
            O => \N__20584\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__2018\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20578\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__20578\,
            I => \N__20575\
        );

    \I__2016\ : Span4Mux_s2_h
    port map (
            O => \N__20575\,
            I => \N__20572\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__20572\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__20569\,
            I => \N__20566\
        );

    \I__2013\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20563\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__20563\,
            I => \N__20560\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__20560\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\
        );

    \I__2010\ : InMux
    port map (
            O => \N__20557\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__2009\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20551\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20548\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__20548\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\
        );

    \I__2006\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20541\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20538\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__20541\,
            I => \N__20535\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__20538\,
            I => \N__20532\
        );

    \I__2002\ : Odrv12
    port map (
            O => \N__20535\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__20532\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8\
        );

    \I__2000\ : InMux
    port map (
            O => \N__20527\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__20524\,
            I => \N__20521\
        );

    \I__1998\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20518\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__20518\,
            I => \N__20515\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__20515\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\
        );

    \I__1995\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20509\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__20509\,
            I => \N__20505\
        );

    \I__1993\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20502\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__20505\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__20502\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8\
        );

    \I__1990\ : InMux
    port map (
            O => \N__20497\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__1989\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20491\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__20491\,
            I => \N__20488\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__20488\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20485\,
            I => \bfn_2_14_0_\
        );

    \I__1985\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20479\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__20476\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\
        );

    \I__1982\ : InMux
    port map (
            O => \N__20473\,
            I => \N__20470\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20467\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__20467\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\
        );

    \I__1979\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20461\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__20461\,
            I => \N__20458\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__20458\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\
        );

    \I__1976\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20452\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20449\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__20449\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\
        );

    \I__1973\ : InMux
    port map (
            O => \N__20446\,
            I => \N__20442\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20445\,
            I => \N__20439\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__20442\,
            I => \N__20436\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__20439\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__20436\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__1968\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20428\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__20428\,
            I => \N__20425\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__20425\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__20422\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12_cascade_\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__20419\,
            I => \N__20416\
        );

    \I__1963\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20412\
        );

    \I__1962\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20409\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__20412\,
            I => \N__20406\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__20409\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__20406\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__1958\ : InMux
    port map (
            O => \N__20401\,
            I => \N__20398\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__20395\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__20392\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13_cascade_\
        );

    \I__1954\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20385\
        );

    \I__1953\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20382\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__20385\,
            I => \N__20379\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__20382\,
            I => \N__20376\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__20379\,
            I => \N__20371\
        );

    \I__1949\ : Span4Mux_v
    port map (
            O => \N__20376\,
            I => \N__20371\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__20371\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__1947\ : InMux
    port map (
            O => \N__20368\,
            I => \N__20365\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__20365\,
            I => \N__20362\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__20362\,
            I => \N__20359\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__20359\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1943\ : InMux
    port map (
            O => \N__20356\,
            I => \N__20350\
        );

    \I__1942\ : InMux
    port map (
            O => \N__20355\,
            I => \N__20350\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__20350\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__1940\ : InMux
    port map (
            O => \N__20347\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__1939\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20341\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__20341\,
            I => \N__20338\
        );

    \I__1937\ : Span4Mux_h
    port map (
            O => \N__20338\,
            I => \N__20335\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__20335\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1935\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20326\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20326\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__20326\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__1932\ : InMux
    port map (
            O => \N__20323\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__1931\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20317\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20314\
        );

    \I__1929\ : Span4Mux_h
    port map (
            O => \N__20314\,
            I => \N__20311\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__20311\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1927\ : InMux
    port map (
            O => \N__20308\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__1926\ : InMux
    port map (
            O => \N__20305\,
            I => \N__20302\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__20302\,
            I => \N__20299\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__20299\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__1923\ : InMux
    port map (
            O => \N__20296\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__1922\ : InMux
    port map (
            O => \N__20293\,
            I => \N__20289\
        );

    \I__1921\ : InMux
    port map (
            O => \N__20292\,
            I => \N__20286\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__20289\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__20286\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__1918\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20275\
        );

    \I__1917\ : InMux
    port map (
            O => \N__20280\,
            I => \N__20275\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__20275\,
            I => \N__20272\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__20272\,
            I => \N__20269\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__20269\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1913\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20263\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__20263\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__20260\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10_cascade_\
        );

    \I__1910\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20253\
        );

    \I__1909\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20250\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__20253\,
            I => \N__20247\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__20250\,
            I => pwm_duty_input_1
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__20247\,
            I => pwm_duty_input_1
        );

    \I__1905\ : InMux
    port map (
            O => \N__20242\,
            I => \N__20239\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__20239\,
            I => \N__20235\
        );

    \I__1903\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20232\
        );

    \I__1902\ : Span4Mux_s1_h
    port map (
            O => \N__20235\,
            I => \N__20229\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__20232\,
            I => pwm_duty_input_0
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__20229\,
            I => pwm_duty_input_0
        );

    \I__1899\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20221\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__20221\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__1897\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20213\
        );

    \I__1896\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20208\
        );

    \I__1895\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20208\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__20213\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__20208\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__1892\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20200\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__20200\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__1890\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20193\
        );

    \I__1889\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20189\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20186\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20183\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__20189\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__20186\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__20183\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__1883\ : InMux
    port map (
            O => \N__20176\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__1882\ : InMux
    port map (
            O => \N__20173\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__1881\ : InMux
    port map (
            O => \N__20170\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__1880\ : InMux
    port map (
            O => \N__20167\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__1879\ : InMux
    port map (
            O => \N__20164\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__1878\ : InMux
    port map (
            O => \N__20161\,
            I => \bfn_2_10_0_\
        );

    \I__1877\ : InMux
    port map (
            O => \N__20158\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__1876\ : InMux
    port map (
            O => \N__20155\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__1875\ : InMux
    port map (
            O => \N__20152\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__1874\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20146\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__20146\,
            I => \N__20143\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__20143\,
            I => \N__20140\
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__20140\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1870\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20134\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__20134\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__1868\ : InMux
    port map (
            O => \N__20131\,
            I => \N__20128\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__20128\,
            I => \N__20125\
        );

    \I__1866\ : Span4Mux_h
    port map (
            O => \N__20125\,
            I => \N__20122\
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__20122\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1864\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20116\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__20116\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__1862\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20110\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__20110\,
            I => \N__20107\
        );

    \I__1860\ : Span4Mux_h
    port map (
            O => \N__20107\,
            I => \N__20104\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__20104\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1858\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20098\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__20098\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__1856\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20092\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__20092\,
            I => \N__20089\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__20089\,
            I => \N__20086\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__20086\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1852\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20080\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__20080\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__1850\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20074\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__20074\,
            I => \N__20071\
        );

    \I__1848\ : Span4Mux_h
    port map (
            O => \N__20071\,
            I => \N__20068\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__20068\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1846\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20062\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__20062\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__1844\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20056\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__20056\,
            I => \N__20053\
        );

    \I__1842\ : Span4Mux_h
    port map (
            O => \N__20053\,
            I => \N__20050\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__20050\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1840\ : InMux
    port map (
            O => \N__20047\,
            I => \N__20044\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__20044\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__1838\ : InMux
    port map (
            O => \N__20041\,
            I => \N__20038\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__20038\,
            I => \N__20035\
        );

    \I__1836\ : Span4Mux_h
    port map (
            O => \N__20035\,
            I => \N__20032\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__20032\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1834\ : InMux
    port map (
            O => \N__20029\,
            I => \N__20026\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__20026\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__1832\ : InMux
    port map (
            O => \N__20023\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__1831\ : InMux
    port map (
            O => \N__20020\,
            I => \bfn_2_6_0_\
        );

    \I__1830\ : InMux
    port map (
            O => \N__20017\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__20014\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__20011\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__1827\ : InMux
    port map (
            O => \N__20008\,
            I => \N__19990\
        );

    \I__1826\ : InMux
    port map (
            O => \N__20007\,
            I => \N__19990\
        );

    \I__1825\ : InMux
    port map (
            O => \N__20006\,
            I => \N__19990\
        );

    \I__1824\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19990\
        );

    \I__1823\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19981\
        );

    \I__1822\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19981\
        );

    \I__1821\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19981\
        );

    \I__1820\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19981\
        );

    \I__1819\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19976\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19976\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__19990\,
            I => \N__19971\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__19981\,
            I => \N__19971\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__19976\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__19971\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__1813\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19963\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__19963\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__1811\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19957\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__19957\,
            I => \N__19954\
        );

    \I__1809\ : Span4Mux_h
    port map (
            O => \N__19954\,
            I => \N__19951\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__19951\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1807\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19945\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__19945\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19939\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__19939\,
            I => \N__19936\
        );

    \I__1803\ : Span4Mux_h
    port map (
            O => \N__19936\,
            I => \N__19933\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__19933\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19927\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__19927\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__1799\ : InMux
    port map (
            O => \N__19924\,
            I => \N__19921\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__19921\,
            I => \N__19918\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__19918\,
            I => \N__19915\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__19915\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19912\,
            I => \N__19909\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__19909\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__1793\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19903\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__19903\,
            I => un7_start_stop_0_a2
        );

    \I__1791\ : InMux
    port map (
            O => \N__19900\,
            I => \bfn_2_5_0_\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19897\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__1789\ : InMux
    port map (
            O => \N__19894\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__1788\ : InMux
    port map (
            O => \N__19891\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__1787\ : InMux
    port map (
            O => \N__19888\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__1786\ : InMux
    port map (
            O => \N__19885\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__1785\ : InMux
    port map (
            O => \N__19882\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__1784\ : InMux
    port map (
            O => \N__19879\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19873\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__19873\,
            I => \N__19870\
        );

    \I__1781\ : Span4Mux_v
    port map (
            O => \N__19870\,
            I => \N__19867\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__19867\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19864\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19861\,
            I => \N__19858\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__19858\,
            I => \N__19855\
        );

    \I__1776\ : Span4Mux_v
    port map (
            O => \N__19855\,
            I => \N__19852\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__19852\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__1774\ : InMux
    port map (
            O => \N__19849\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19846\,
            I => \N__19843\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19843\,
            I => \N__19840\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__19840\,
            I => \N__19837\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__19837\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19834\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__1768\ : InMux
    port map (
            O => \N__19831\,
            I => \N__19828\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__19828\,
            I => \N__19825\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__19825\,
            I => \N__19822\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__19822\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__1764\ : InMux
    port map (
            O => \N__19819\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__19816\,
            I => \N__19813\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19810\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__19810\,
            I => \N__19807\
        );

    \I__1760\ : Span12Mux_v
    port map (
            O => \N__19807\,
            I => \N__19804\
        );

    \I__1759\ : Odrv12
    port map (
            O => \N__19804\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19801\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__1757\ : InMux
    port map (
            O => \N__19798\,
            I => \bfn_1_13_0_\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19792\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__19792\,
            I => \N__19789\
        );

    \I__1754\ : Span4Mux_v
    port map (
            O => \N__19789\,
            I => \N__19786\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__19786\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__1752\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19780\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__19780\,
            I => \N__19777\
        );

    \I__1750\ : Span4Mux_v
    port map (
            O => \N__19777\,
            I => \N__19769\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__19776\,
            I => \N__19765\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__19775\,
            I => \N__19762\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__19774\,
            I => \N__19758\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__19773\,
            I => \N__19755\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__19772\,
            I => \N__19752\
        );

    \I__1744\ : Span4Mux_v
    port map (
            O => \N__19769\,
            I => \N__19749\
        );

    \I__1743\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19746\
        );

    \I__1742\ : InMux
    port map (
            O => \N__19765\,
            I => \N__19741\
        );

    \I__1741\ : InMux
    port map (
            O => \N__19762\,
            I => \N__19741\
        );

    \I__1740\ : InMux
    port map (
            O => \N__19761\,
            I => \N__19732\
        );

    \I__1739\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19732\
        );

    \I__1738\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19732\
        );

    \I__1737\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19732\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__19749\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__19746\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__19741\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__19732\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__19723\,
            I => \N__19720\
        );

    \I__1731\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19717\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19713\
        );

    \I__1729\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19710\
        );

    \I__1728\ : Span4Mux_v
    port map (
            O => \N__19713\,
            I => \N__19707\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__19710\,
            I => \N__19704\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__19707\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__19704\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__1724\ : InMux
    port map (
            O => \N__19699\,
            I => \N__19696\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__19696\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__1722\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19690\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__19690\,
            I => \N_42_i_i\
        );

    \I__1720\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19684\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19681\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__19681\,
            I => \N__19678\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__19678\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__19675\,
            I => \N__19672\
        );

    \I__1715\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19669\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__19669\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__1713\ : InMux
    port map (
            O => \N__19666\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__1712\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19660\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__19660\,
            I => \N__19657\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__19657\,
            I => \N__19654\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__19654\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__19651\,
            I => \N__19648\
        );

    \I__1707\ : InMux
    port map (
            O => \N__19648\,
            I => \N__19645\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__19645\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__1705\ : InMux
    port map (
            O => \N__19642\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__1704\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19636\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__19636\,
            I => \N__19633\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__19633\,
            I => \N__19630\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__19630\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__19627\,
            I => \N__19624\
        );

    \I__1699\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19621\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__19621\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19618\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__1696\ : InMux
    port map (
            O => \N__19615\,
            I => \N__19612\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__19612\,
            I => \N__19609\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__19609\,
            I => \N__19606\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__19606\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__19603\,
            I => \N__19600\
        );

    \I__1691\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19597\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__19597\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__1689\ : InMux
    port map (
            O => \N__19594\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__1688\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19588\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__19588\,
            I => \N__19585\
        );

    \I__1686\ : Span4Mux_v
    port map (
            O => \N__19585\,
            I => \N__19582\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__19582\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__19579\,
            I => \N__19576\
        );

    \I__1683\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19573\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__19573\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__1681\ : InMux
    port map (
            O => \N__19570\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__1680\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19564\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__19564\,
            I => \N__19561\
        );

    \I__1678\ : Span4Mux_v
    port map (
            O => \N__19561\,
            I => \N__19558\
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__19558\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__19555\,
            I => \N__19552\
        );

    \I__1675\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19549\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__19549\,
            I => \N__19546\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__19546\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__1672\ : InMux
    port map (
            O => \N__19543\,
            I => \bfn_1_12_0_\
        );

    \I__1671\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19537\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__19537\,
            I => \N__19534\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__19534\,
            I => \N__19531\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__19531\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__1666\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19522\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__19522\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19519\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__1663\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19513\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__19513\,
            I => \N__19510\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__19510\,
            I => \N__19507\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__19507\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__1659\ : InMux
    port map (
            O => \N__19504\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__1658\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19498\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__19498\,
            I => \N__19495\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__19495\,
            I => \N__19492\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__19492\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__19489\,
            I => \N__19486\
        );

    \I__1653\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19483\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__19483\,
            I => \N__19480\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__19480\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__1650\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19474\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19471\
        );

    \I__1648\ : Span4Mux_v
    port map (
            O => \N__19471\,
            I => \N__19468\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__19468\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__19465\,
            I => \N__19462\
        );

    \I__1645\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19459\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__19459\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__1643\ : InMux
    port map (
            O => \N__19456\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__1642\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19450\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__19450\,
            I => \N__19447\
        );

    \I__1640\ : Span4Mux_v
    port map (
            O => \N__19447\,
            I => \N__19444\
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__19444\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__19441\,
            I => \N__19438\
        );

    \I__1637\ : InMux
    port map (
            O => \N__19438\,
            I => \N__19435\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__19435\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__1635\ : InMux
    port map (
            O => \N__19432\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__1634\ : IoInMux
    port map (
            O => \N__19429\,
            I => \N__19426\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__19426\,
            I => \N__19423\
        );

    \I__1632\ : Span4Mux_s3_v
    port map (
            O => \N__19423\,
            I => \N__19420\
        );

    \I__1631\ : Span4Mux_h
    port map (
            O => \N__19420\,
            I => \N__19417\
        );

    \I__1630\ : Sp12to4
    port map (
            O => \N__19417\,
            I => \N__19414\
        );

    \I__1629\ : Span12Mux_v
    port map (
            O => \N__19414\,
            I => \N__19411\
        );

    \I__1628\ : Span12Mux_v
    port map (
            O => \N__19411\,
            I => \N__19408\
        );

    \I__1627\ : Odrv12
    port map (
            O => \N__19408\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1626\ : IoInMux
    port map (
            O => \N__19405\,
            I => \N__19402\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__1624\ : IoSpan4Mux
    port map (
            O => \N__19399\,
            I => \N__19396\
        );

    \I__1623\ : IoSpan4Mux
    port map (
            O => \N__19396\,
            I => \N__19393\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__19393\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_10_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_10_25_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_3_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_3_10_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_3_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_7_0_\
        );

    \IN_MUX_bfv_3_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_3_8_0_\
        );

    \IN_MUX_bfv_2_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_5_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_7_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_7_22_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_8_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_8_23_0_\
        );

    \IN_MUX_bfv_8_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_8_24_0_\
        );

    \IN_MUX_bfv_13_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_4_0_\
        );

    \IN_MUX_bfv_13_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            carryinitout => \bfn_13_5_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_12_10_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19429\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19405\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26158\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_397_i_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__34831\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_166_i_g\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__28960\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_399_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__28304\,
            CLKHFEN => \N__28308\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__28315\,
            RGB2PWM => \N__19693\,
            RGB1 => rgb_g_wire,
            CURREN => \N__28309\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__19906\,
            RGB0PWM => \N__49588\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__19783\,
            in1 => \N__19716\,
            in2 => \_gnd_net_\,
            in3 => \N__21378\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23176\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49977\,
            ce => 'H',
            sr => \N__49496\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__23175\,
            in1 => \N__22123\,
            in2 => \N__22578\,
            in3 => \N__22358\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49975\,
            ce => 'H',
            sr => \N__49516\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__21768\,
            in1 => \N__22435\,
            in2 => \N__22182\,
            in3 => \N__22266\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => 'H',
            sr => \N__49520\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__22420\,
            in1 => \N__21769\,
            in2 => \N__22183\,
            in3 => \N__22267\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => 'H',
            sr => \N__49520\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__21253\,
            in1 => \N__22355\,
            in2 => \N__21235\,
            in3 => \N__22696\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => 'H',
            sr => \N__49520\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__23169\,
            in1 => \N__22615\,
            in2 => \N__22359\,
            in3 => \N__22121\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => 'H',
            sr => \N__49520\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__22119\,
            in1 => \N__23168\,
            in2 => \N__22657\,
            in3 => \N__22356\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => 'H',
            sr => \N__49520\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__23170\,
            in1 => \N__22543\,
            in2 => \N__22360\,
            in3 => \N__22122\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => 'H',
            sr => \N__49520\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__22120\,
            in1 => \N__23171\,
            in2 => \N__22507\,
            in3 => \N__22357\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49973\,
            ce => 'H',
            sr => \N__49520\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19501\,
            in2 => \N__19489\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19477\,
            in2 => \N__19465\,
            in3 => \N__19456\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19453\,
            in2 => \N__19441\,
            in3 => \N__19432\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19687\,
            in2 => \N__19675\,
            in3 => \N__19666\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19663\,
            in2 => \N__19651\,
            in3 => \N__19642\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19639\,
            in2 => \N__19627\,
            in3 => \N__19618\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19615\,
            in2 => \N__19603\,
            in3 => \N__19594\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19591\,
            in2 => \N__19579\,
            in3 => \N__19570\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19567\,
            in2 => \N__19555\,
            in3 => \N__19543\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19540\,
            in2 => \N__19528\,
            in3 => \N__19519\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19516\,
            in2 => \N__19772\,
            in3 => \N__19504\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19876\,
            in2 => \N__19775\,
            in3 => \N__19864\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19861\,
            in2 => \N__19773\,
            in3 => \N__19849\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19846\,
            in2 => \N__19776\,
            in3 => \N__19834\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19831\,
            in2 => \N__19774\,
            in3 => \N__19819\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19761\,
            in2 => \N__19816\,
            in3 => \N__19801\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20581\,
            in1 => \N__19699\,
            in2 => \_gnd_net_\,
            in3 => \N__19798\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__19795\,
            in1 => \N__19768\,
            in2 => \N__19723\,
            in3 => \N__21411\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.N_42_i_i_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__33156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49586\,
            lcout => \N_42_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__33160\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49587\,
            lcout => un7_start_stop_0_a2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20005\,
            in1 => \N__20834\,
            in2 => \_gnd_net_\,
            in3 => \N__19900\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_5_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__49978\,
            ce => 'H',
            sr => \N__49483\
        );

    \pwm_generator_inst.counter_1_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20001\,
            in1 => \N__20807\,
            in2 => \_gnd_net_\,
            in3 => \N__19897\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__49978\,
            ce => 'H',
            sr => \N__49483\
        );

    \pwm_generator_inst.counter_2_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20006\,
            in1 => \N__20762\,
            in2 => \_gnd_net_\,
            in3 => \N__19894\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__49978\,
            ce => 'H',
            sr => \N__49483\
        );

    \pwm_generator_inst.counter_3_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20002\,
            in1 => \N__20738\,
            in2 => \_gnd_net_\,
            in3 => \N__19891\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__49978\,
            ce => 'H',
            sr => \N__49483\
        );

    \pwm_generator_inst.counter_4_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20007\,
            in1 => \N__20699\,
            in2 => \_gnd_net_\,
            in3 => \N__19888\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__49978\,
            ce => 'H',
            sr => \N__49483\
        );

    \pwm_generator_inst.counter_5_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20003\,
            in1 => \N__20672\,
            in2 => \_gnd_net_\,
            in3 => \N__19885\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__49978\,
            ce => 'H',
            sr => \N__49483\
        );

    \pwm_generator_inst.counter_6_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20008\,
            in1 => \N__21011\,
            in2 => \_gnd_net_\,
            in3 => \N__19882\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__49978\,
            ce => 'H',
            sr => \N__49483\
        );

    \pwm_generator_inst.counter_7_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20004\,
            in1 => \N__20984\,
            in2 => \_gnd_net_\,
            in3 => \N__19879\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__49978\,
            ce => 'H',
            sr => \N__49483\
        );

    \pwm_generator_inst.counter_8_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20000\,
            in1 => \N__20952\,
            in2 => \_gnd_net_\,
            in3 => \N__20020\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__49976\,
            ce => 'H',
            sr => \N__49490\
        );

    \pwm_generator_inst.counter_9_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__20925\,
            in1 => \N__19999\,
            in2 => \_gnd_net_\,
            in3 => \N__20017\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49976\,
            ce => 'H',
            sr => \N__49490\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20838\,
            in2 => \_gnd_net_\,
            in3 => \N__20770\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__20701\,
            in1 => \N__20740\,
            in2 => \N__20014\,
            in3 => \N__20809\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19966\,
            in1 => \N__21013\,
            in2 => \N__20011\,
            in3 => \N__20674\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20985\,
            in1 => \N__20921\,
            in2 => \_gnd_net_\,
            in3 => \N__20948\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19948\,
            in2 => \_gnd_net_\,
            in3 => \N__19960\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19930\,
            in2 => \_gnd_net_\,
            in3 => \N__19942\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19912\,
            in2 => \_gnd_net_\,
            in3 => \N__19924\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20149\,
            in1 => \N__20137\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20119\,
            in2 => \_gnd_net_\,
            in3 => \N__20131\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20101\,
            in2 => \_gnd_net_\,
            in3 => \N__20113\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20083\,
            in2 => \_gnd_net_\,
            in3 => \N__20095\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20065\,
            in2 => \_gnd_net_\,
            in3 => \N__20077\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20047\,
            in2 => \_gnd_net_\,
            in3 => \N__20059\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20029\,
            in2 => \_gnd_net_\,
            in3 => \N__20041\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20292\,
            in2 => \_gnd_net_\,
            in3 => \N__20023\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__21998\,
            in1 => \N__20389\,
            in2 => \_gnd_net_\,
            in3 => \N__20176\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20446\,
            in2 => \_gnd_net_\,
            in3 => \N__20173\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20419\,
            in3 => \N__20170\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21204\,
            in2 => \_gnd_net_\,
            in3 => \N__20167\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22059\,
            in2 => \_gnd_net_\,
            in3 => \N__20164\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21041\,
            in2 => \_gnd_net_\,
            in3 => \N__20161\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20216\,
            in2 => \_gnd_net_\,
            in3 => \N__20158\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20197\,
            in2 => \_gnd_net_\,
            in3 => \N__20155\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20152\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20280\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20281\,
            in1 => \N__20266\,
            in2 => \N__20260\,
            in3 => \N__21981\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__21744\,
            in1 => \N__20256\,
            in2 => \_gnd_net_\,
            in3 => \N__20238\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__20224\,
            in1 => \N__20217\,
            in2 => \N__22003\,
            in3 => \N__20545\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20218\,
            in2 => \_gnd_net_\,
            in3 => \N__20544\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__20192\,
            in1 => \N__20512\,
            in2 => \N__22004\,
            in3 => \N__20203\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21063\,
            in2 => \_gnd_net_\,
            in3 => \N__21045\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20196\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__22058\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22026\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20355\,
            in2 => \_gnd_net_\,
            in3 => \N__20445\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20356\,
            in1 => \N__20431\,
            in2 => \N__20422\,
            in3 => \N__21967\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20331\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20332\,
            in1 => \N__20401\,
            in2 => \N__20392\,
            in3 => \N__21968\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20388\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20368\,
            in2 => \_gnd_net_\,
            in3 => \N__20347\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20344\,
            in2 => \_gnd_net_\,
            in3 => \N__20323\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20320\,
            in2 => \_gnd_net_\,
            in3 => \N__20308\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20305\,
            in2 => \_gnd_net_\,
            in3 => \N__20296\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28277\,
            in2 => \N__20569\,
            in3 => \N__20557\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20554\,
            in2 => \N__28310\,
            in3 => \N__20527\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28281\,
            in2 => \N__20524\,
            in3 => \N__20497\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20494\,
            in2 => \_gnd_net_\,
            in3 => \N__20485\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20482\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20473\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20464\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20455\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20647\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20638\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20629\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20620\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20611\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20602\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20593\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20584\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__21598\,
            in1 => \N__20851\,
            in2 => \N__21428\,
            in3 => \N__21813\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__21599\,
            in1 => \N__21124\,
            in2 => \N__21429\,
            in3 => \N__21814\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20815\,
            in2 => \N__21145\,
            in3 => \N__20839\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_3_7_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20788\,
            in2 => \N__21472\,
            in3 => \N__20808\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20746\,
            in2 => \N__20782\,
            in3 => \N__20769\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20739\,
            in1 => \N__20707\,
            in2 => \N__20719\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20700\,
            in1 => \N__20680\,
            in2 => \N__21487\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20673\,
            in1 => \N__20653\,
            in2 => \N__21523\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21012\,
            in1 => \N__20992\,
            in2 => \N__21508\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21277\,
            in2 => \N__20962\,
            in3 => \N__20986\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20953\,
            in1 => \N__20932\,
            in2 => \N__21448\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_3_8_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20905\,
            in2 => \N__21544\,
            in3 => \N__20926\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20899\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49974\,
            ce => 'H',
            sr => \N__49497\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20875\,
            in2 => \N__22013\,
            in3 => \N__22005\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20869\,
            in2 => \_gnd_net_\,
            in3 => \N__20863\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20860\,
            in2 => \_gnd_net_\,
            in3 => \N__20842\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21136\,
            in2 => \_gnd_net_\,
            in3 => \N__21115\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21259\,
            in2 => \_gnd_net_\,
            in3 => \N__21112\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21922\,
            in2 => \_gnd_net_\,
            in3 => \N__21109\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21019\,
            in2 => \_gnd_net_\,
            in3 => \N__21106\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21103\,
            in2 => \_gnd_net_\,
            in3 => \N__21097\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21094\,
            in2 => \_gnd_net_\,
            in3 => \N__21088\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271\,
            ltout => OPEN,
            carryin => \bfn_3_10_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__21085\,
            in1 => \N__21079\,
            in2 => \N__22015\,
            in3 => \N__21067\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22608\,
            in1 => \N__22502\,
            in2 => \N__22579\,
            in3 => \N__21271\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__21064\,
            in1 => \N__22009\,
            in2 => \N__21046\,
            in3 => \N__21025\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__22650\,
            in1 => \N__22524\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__21840\,
            in1 => \N__21915\,
            in2 => \N__21879\,
            in3 => \N__21661\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__21265\,
            in1 => \N__21220\,
            in2 => \N__22014\,
            in3 => \N__21205\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__23165\,
            in1 => \N__21246\,
            in2 => \N__22240\,
            in3 => \N__22329\,
            lcout => \current_shift_inst.PI_CTRL.N_153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__23167\,
            in1 => \N__22692\,
            in2 => \N__22230\,
            in3 => \N__22096\,
            lcout => \current_shift_inst.PI_CTRL.N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__23166\,
            in1 => \_gnd_net_\,
            in2 => \N__22231\,
            in3 => \N__22095\,
            lcout => \current_shift_inst.PI_CTRL.N_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__21197\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21216\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21181\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__21600\,
            in1 => \N__21154\,
            in2 => \N__21433\,
            in3 => \N__21807\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__21806\,
            in1 => \N__21607\,
            in2 => \N__21556\,
            in3 => \N__21423\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__21802\,
            in1 => \N__21603\,
            in2 => \N__21532\,
            in3 => \N__21419\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__21604\,
            in1 => \N__21514\,
            in2 => \N__21431\,
            in3 => \N__21803\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__21801\,
            in1 => \N__21602\,
            in2 => \N__21496\,
            in3 => \N__21418\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__21601\,
            in1 => \N__21478\,
            in2 => \N__21430\,
            in3 => \N__21800\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110011"
        )
    port map (
            in0 => \N__21805\,
            in1 => \N__21606\,
            in2 => \N__21463\,
            in3 => \N__21424\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__21605\,
            in1 => \N__21439\,
            in2 => \N__21432\,
            in3 => \N__21804\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__22189\,
            in1 => \N__22607\,
            in2 => \N__22542\,
            in3 => \N__22571\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__22072\,
            in1 => \N__22063\,
            in2 => \N__22036\,
            in3 => \N__21999\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21916\,
            in1 => \N__21880\,
            in2 => \N__21727\,
            in3 => \N__21844\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__21691\,
            in1 => \N__22383\,
            in2 => \N__21817\,
            in3 => \N__21648\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__22257\,
            in1 => \N__21761\,
            in2 => \N__22174\,
            in3 => \N__22405\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49967\,
            ce => 'H',
            sr => \N__49506\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__21723\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21686\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101011"
        )
    port map (
            in0 => \N__21655\,
            in1 => \N__22382\,
            in2 => \N__21649\,
            in3 => \N__21616\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22777\,
            in2 => \_gnd_net_\,
            in3 => \N__22800\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22941\,
            in1 => \N__22288\,
            in2 => \N__21562\,
            in3 => \N__22918\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22300\,
            in1 => \N__22282\,
            in2 => \N__21559\,
            in3 => \N__22246\,
            lcout => \current_shift_inst.PI_CTRL.N_53\,
            ltout => \current_shift_inst.PI_CTRL.N_53_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000100"
        )
    port map (
            in0 => \N__22725\,
            in1 => \N__22156\,
            in2 => \N__22270\,
            in3 => \N__22138\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23052\,
            in1 => \N__22447\,
            in2 => \N__23074\,
            in3 => \N__23245\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22690\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22724\,
            lcout => \current_shift_inst.PI_CTRL.N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__22223\,
            in1 => \N__23142\,
            in2 => \_gnd_net_\,
            in3 => \N__22691\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26207\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__49521\
        );

    \delay_measurement_inst.start_timer_hc_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26206\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22207\,
            ce => 'H',
            sr => \N__49521\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22198\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49972\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22503\,
            in2 => \_gnd_net_\,
            in3 => \N__22640\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101010001"
        )
    port map (
            in0 => \N__22175\,
            in1 => \N__22137\,
            in2 => \N__22118\,
            in3 => \N__22726\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49962\,
            ce => 'H',
            sr => \N__49498\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23244\,
            in1 => \N__22306\,
            in2 => \N__22942\,
            in3 => \N__22294\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22276\,
            in1 => \N__22312\,
            in2 => \N__22363\,
            in3 => \N__22453\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23094\,
            in1 => \N__22872\,
            in2 => \N__22896\,
            in3 => \N__22746\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23013\,
            in1 => \N__23028\,
            in2 => \N__23221\,
            in3 => \N__23070\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23029\,
            in1 => \N__22873\,
            in2 => \N__22897\,
            in3 => \N__23014\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22917\,
            in2 => \_gnd_net_\,
            in3 => \N__22470\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22471\,
            in1 => \N__22824\,
            in2 => \N__22855\,
            in3 => \N__23220\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22996\,
            in1 => \N__23098\,
            in2 => \N__22981\,
            in3 => \N__22750\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23194\,
            in1 => \N__22776\,
            in2 => \N__22960\,
            in3 => \N__22801\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22995\,
            in1 => \N__23053\,
            in2 => \N__22980\,
            in3 => \N__22441\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23193\,
            in2 => \_gnd_net_\,
            in3 => \N__22959\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22825\,
            in2 => \_gnd_net_\,
            in3 => \N__22851\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__37664\,
            in1 => \N__37285\,
            in2 => \_gnd_net_\,
            in3 => \N__26689\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49970\,
            ce => 'H',
            sr => \N__49452\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29841\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30312\,
            in1 => \N__35456\,
            in2 => \N__33813\,
            in3 => \N__29714\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25411\,
            in2 => \N__24577\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__49957\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25402\,
            in2 => \N__29434\,
            in3 => \N__22408\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__49957\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29257\,
            in2 => \N__25423\,
            in3 => \N__22393\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__49957\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23407\,
            in2 => \N__34801\,
            in3 => \N__22699\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__49957\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23413\,
            in2 => \N__29587\,
            in3 => \N__22660\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__49957\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23395\,
            in2 => \N__29641\,
            in3 => \N__22618\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__49957\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23419\,
            in2 => \N__29347\,
            in3 => \N__22582\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__49957\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23401\,
            in2 => \N__33955\,
            in3 => \N__22546\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__49957\,
            ce => 'H',
            sr => \N__49474\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25459\,
            in2 => \N__37114\,
            in3 => \N__22510\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__49951\,
            ce => 'H',
            sr => \N__49484\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24640\,
            in2 => \N__38110\,
            in3 => \N__22474\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__49951\,
            ce => 'H',
            sr => \N__49484\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24667\,
            in2 => \N__33871\,
            in3 => \N__22456\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__49951\,
            ce => 'H',
            sr => \N__49484\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24649\,
            in2 => \N__35284\,
            in3 => \N__22921\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__49951\,
            ce => 'H',
            sr => \N__49484\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25393\,
            in2 => \N__29797\,
            in3 => \N__22900\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__49951\,
            ce => 'H',
            sr => \N__49484\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24658\,
            in2 => \N__38179\,
            in3 => \N__22876\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__49951\,
            ce => 'H',
            sr => \N__49484\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25480\,
            in2 => \N__29215\,
            in3 => \N__22858\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__49951\,
            ce => 'H',
            sr => \N__49484\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29490\,
            in2 => \N__25518\,
            in3 => \N__22828\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__49951\,
            ce => 'H',
            sr => \N__49484\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25519\,
            in2 => \N__38041\,
            in3 => \N__22804\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33718\,
            in2 => \N__25551\,
            in3 => \N__22780\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25523\,
            in2 => \N__35130\,
            in3 => \N__22753\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35655\,
            in2 => \N__25552\,
            in3 => \N__22729\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25527\,
            in2 => \N__34015\,
            in3 => \N__23077\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33817\,
            in2 => \N__25553\,
            in3 => \N__23056\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25531\,
            in2 => \N__29857\,
            in3 => \N__23032\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30003\,
            in2 => \N__25554\,
            in3 => \N__23017\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__49947\,
            ce => 'H',
            sr => \N__49491\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35457\,
            in2 => \N__25555\,
            in3 => \N__22999\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__49943\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25538\,
            in2 => \N__30316\,
            in3 => \N__22984\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__49943\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29718\,
            in2 => \N__25556\,
            in3 => \N__22963\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__49943\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25542\,
            in2 => \N__34090\,
            in3 => \N__22945\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__49943\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27148\,
            in2 => \N__25557\,
            in3 => \N__23224\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__49943\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25546\,
            in2 => \N__27193\,
            in3 => \N__23197\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__49943\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25384\,
            in2 => \N__25558\,
            in3 => \N__23182\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__49943\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37500\,
            in1 => \N__25550\,
            in2 => \_gnd_net_\,
            in3 => \N__23179\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => 'H',
            sr => \N__49499\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30745\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24756\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25922\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30829\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27334\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24802\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__31985\,
            in1 => \N__24834\,
            in2 => \N__27436\,
            in3 => \N__24813\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23890\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49931\,
            ce => \N__27634\,
            sr => \N__49509\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__31986\,
            in1 => \N__26415\,
            in2 => \N__28000\,
            in3 => \N__32667\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30919\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30512\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31351\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25958\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26302\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26065\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31642\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32146\,
            in1 => \N__26474\,
            in2 => \N__32726\,
            in3 => \N__26438\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31048\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32141\,
            in1 => \N__31169\,
            in2 => \N__32725\,
            in3 => \N__31130\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__30490\,
            in1 => \N__32140\,
            in2 => \N__32728\,
            in3 => \N__30513\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__25826\,
            in1 => \N__32711\,
            in2 => \N__32155\,
            in3 => \N__25790\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27266\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32142\,
            in1 => \N__26376\,
            in2 => \N__32727\,
            in3 => \N__26330\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24884\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24942\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31168\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25825\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26368\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31781\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31543\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26473\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24704\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23914\,
            in2 => \N__23862\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__49903\,
            ce => \N__27631\,
            sr => \N__49528\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23886\,
            in2 => \N__23835\,
            in3 => \N__23248\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__49903\,
            ce => \N__27631\,
            sr => \N__49528\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23805\,
            in2 => \N__23863\,
            in3 => \N__23275\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__49903\,
            ce => \N__27631\,
            sr => \N__49528\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23778\,
            in2 => \N__23836\,
            in3 => \N__23272\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__49903\,
            ce => \N__27631\,
            sr => \N__49528\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23751\,
            in2 => \N__23809\,
            in3 => \N__23269\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__49903\,
            ce => \N__27631\,
            sr => \N__49528\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24123\,
            in2 => \N__23782\,
            in3 => \N__23266\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__49903\,
            ce => \N__27631\,
            sr => \N__49528\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24099\,
            in2 => \N__23755\,
            in3 => \N__23263\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__49903\,
            ce => \N__27631\,
            sr => \N__49528\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24124\,
            in2 => \N__24076\,
            in3 => \N__23260\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__49903\,
            ce => \N__27631\,
            sr => \N__49528\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24042\,
            in2 => \N__24103\,
            in3 => \N__23257\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__49898\,
            ce => \N__27630\,
            sr => \N__49533\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24018\,
            in2 => \N__24075\,
            in3 => \N__23254\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__49898\,
            ce => \N__27630\,
            sr => \N__49533\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24043\,
            in2 => \N__23995\,
            in3 => \N__23251\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__49898\,
            ce => \N__27630\,
            sr => \N__49533\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23964\,
            in2 => \N__24022\,
            in3 => \N__23302\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__49898\,
            ce => \N__27630\,
            sr => \N__49533\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23994\,
            in2 => \N__23940\,
            in3 => \N__23299\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__49898\,
            ce => \N__27630\,
            sr => \N__49533\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24351\,
            in2 => \N__23968\,
            in3 => \N__23296\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__49898\,
            ce => \N__27630\,
            sr => \N__49533\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24327\,
            in2 => \N__23941\,
            in3 => \N__23293\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__49898\,
            ce => \N__27630\,
            sr => \N__49533\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24352\,
            in2 => \N__24303\,
            in3 => \N__23290\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__49898\,
            ce => \N__27630\,
            sr => \N__49533\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24273\,
            in2 => \N__24331\,
            in3 => \N__23287\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__49892\,
            ce => \N__27628\,
            sr => \N__49537\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24249\,
            in2 => \N__24304\,
            in3 => \N__23284\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__49892\,
            ce => \N__27628\,
            sr => \N__49537\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24274\,
            in2 => \N__24226\,
            in3 => \N__23281\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__49892\,
            ce => \N__27628\,
            sr => \N__49537\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24195\,
            in2 => \N__24253\,
            in3 => \N__23278\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__49892\,
            ce => \N__27628\,
            sr => \N__49537\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24225\,
            in2 => \N__24171\,
            in3 => \N__23329\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__49892\,
            ce => \N__27628\,
            sr => \N__49537\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24144\,
            in2 => \N__24199\,
            in3 => \N__23326\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__49892\,
            ce => \N__27628\,
            sr => \N__49537\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24504\,
            in2 => \N__24172\,
            in3 => \N__23323\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__49892\,
            ce => \N__27628\,
            sr => \N__49537\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24145\,
            in2 => \N__24480\,
            in3 => \N__23320\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__49892\,
            ce => \N__27628\,
            sr => \N__49537\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24450\,
            in2 => \N__24508\,
            in3 => \N__23317\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_7_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__49885\,
            ce => \N__27627\,
            sr => \N__49541\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24426\,
            in2 => \N__24481\,
            in3 => \N__23314\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__49885\,
            ce => \N__27627\,
            sr => \N__49541\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24451\,
            in2 => \N__24403\,
            in3 => \N__23311\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__49885\,
            ce => \N__27627\,
            sr => \N__49541\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24379\,
            in2 => \N__24430\,
            in3 => \N__23308\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__49885\,
            ce => \N__27627\,
            sr => \N__49541\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23305\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23380\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49971\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__37663\,
            in1 => \N__37234\,
            in2 => \_gnd_net_\,
            in3 => \N__26728\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49968\,
            ce => 'H',
            sr => \N__49444\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38037\,
            in1 => \N__29204\,
            in2 => \N__38174\,
            in3 => \N__29997\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27147\,
            in1 => \N__23365\,
            in2 => \N__23368\,
            in3 => \N__34084\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25380\,
            in2 => \_gnd_net_\,
            in3 => \N__29793\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23359\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49958\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37488\,
            in1 => \N__35123\,
            in2 => \N__29852\,
            in3 => \N__35656\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23347\,
            in1 => \N__23341\,
            in2 => \N__23335\,
            in3 => \N__23425\,
            lcout => \current_shift_inst.PI_CTRL.N_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37107\,
            in1 => \N__33936\,
            in2 => \N__29346\,
            in3 => \N__38103\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__29582\,
            in1 => \N__34796\,
            in2 => \N__23332\,
            in3 => \N__29637\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33862\,
            in1 => \N__24607\,
            in2 => \N__23428\,
            in3 => \N__27185\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30148\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49467\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29916\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49467\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33231\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49467\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30119\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49467\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29886\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49467\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27485\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__27486\,
            in1 => \_gnd_net_\,
            in2 => \N__23389\,
            in3 => \N__30656\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23386\,
            in2 => \N__27527\,
            in3 => \N__27528\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23725\,
            in2 => \_gnd_net_\,
            in3 => \N__23494\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23491\,
            in2 => \_gnd_net_\,
            in3 => \N__23485\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23482\,
            in2 => \_gnd_net_\,
            in3 => \N__23476\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23473\,
            in2 => \_gnd_net_\,
            in3 => \N__23467\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23464\,
            in2 => \_gnd_net_\,
            in3 => \N__23452\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23449\,
            in2 => \_gnd_net_\,
            in3 => \N__23443\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23440\,
            in2 => \_gnd_net_\,
            in3 => \N__23434\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23686\,
            in2 => \_gnd_net_\,
            in3 => \N__23431\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23701\,
            in3 => \N__23563\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23560\,
            in2 => \_gnd_net_\,
            in3 => \N__23554\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23713\,
            in2 => \_gnd_net_\,
            in3 => \N__23551\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23548\,
            in2 => \_gnd_net_\,
            in3 => \N__23542\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23539\,
            in2 => \_gnd_net_\,
            in3 => \N__23533\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23530\,
            in2 => \_gnd_net_\,
            in3 => \N__23524\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23521\,
            in2 => \_gnd_net_\,
            in3 => \N__23515\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23512\,
            in2 => \_gnd_net_\,
            in3 => \N__23506\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23503\,
            in2 => \_gnd_net_\,
            in3 => \N__23497\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23641\,
            in2 => \_gnd_net_\,
            in3 => \N__23632\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23629\,
            in2 => \_gnd_net_\,
            in3 => \N__23620\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23617\,
            in2 => \_gnd_net_\,
            in3 => \N__23608\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25843\,
            in2 => \_gnd_net_\,
            in3 => \N__23605\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23602\,
            in2 => \_gnd_net_\,
            in3 => \N__23593\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23590\,
            in2 => \_gnd_net_\,
            in3 => \N__23584\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23581\,
            in2 => \_gnd_net_\,
            in3 => \N__23575\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23572\,
            in2 => \_gnd_net_\,
            in3 => \N__23566\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23677\,
            in2 => \_gnd_net_\,
            in3 => \N__23671\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23668\,
            in2 => \_gnd_net_\,
            in3 => \N__23662\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23659\,
            in2 => \_gnd_net_\,
            in3 => \N__23650\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23647\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23644\,
            in3 => \N__32138\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30620\,
            in1 => \N__30749\,
            in2 => \_gnd_net_\,
            in3 => \N__30714\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__30619\,
            in1 => \N__25995\,
            in2 => \_gnd_net_\,
            in3 => \N__25952\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__27335\,
            in1 => \N__30616\,
            in2 => \_gnd_net_\,
            in3 => \N__27303\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32108\,
            in1 => \N__27267\,
            in2 => \_gnd_net_\,
            in3 => \N__27225\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__25871\,
            in1 => \N__30618\,
            in2 => \_gnd_net_\,
            in3 => \N__25915\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30615\,
            in1 => \N__30830\,
            in2 => \_gnd_net_\,
            in3 => \N__30798\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30622\,
            in1 => \N__31406\,
            in2 => \_gnd_net_\,
            in3 => \N__31449\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30617\,
            in1 => \N__24711\,
            in2 => \_gnd_net_\,
            in3 => \N__24687\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30621\,
            in1 => \N__24752\,
            in2 => \_gnd_net_\,
            in3 => \N__24787\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__30923\,
            in1 => \N__30643\,
            in2 => \_gnd_net_\,
            in3 => \N__30888\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30645\,
            in1 => \N__31059\,
            in2 => \_gnd_net_\,
            in3 => \N__31088\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30981\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__30647\,
            in1 => \_gnd_net_\,
            in2 => \N__31788\,
            in3 => \N__31829\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__26066\,
            in1 => \N__30646\,
            in2 => \_gnd_net_\,
            in3 => \N__26028\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30648\,
            in1 => \N__31228\,
            in2 => \_gnd_net_\,
            in3 => \N__31266\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__27558\,
            in1 => \N__30642\,
            in2 => \_gnd_net_\,
            in3 => \N__27599\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30644\,
            in1 => \N__26303\,
            in2 => \_gnd_net_\,
            in3 => \N__26258\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__31653\,
            in1 => \N__31595\,
            in2 => \_gnd_net_\,
            in3 => \N__30655\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27557\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26112\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30654\,
            in1 => \N__31544\,
            in2 => \_gnd_net_\,
            in3 => \N__31512\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32156\,
            in1 => \N__26369\,
            in2 => \_gnd_net_\,
            in3 => \N__26337\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31396\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__32158\,
            in1 => \_gnd_net_\,
            in2 => \N__26481\,
            in3 => \N__26442\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__25827\,
            in1 => \N__32157\,
            in2 => \_gnd_net_\,
            in3 => \N__25794\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23913\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49893\,
            ce => \N__27629\,
            sr => \N__49529\
        );

    \current_shift_inst.timer_s1.counter_0_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25325\,
            in1 => \N__23912\,
            in2 => \_gnd_net_\,
            in3 => \N__23893\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__49886\,
            ce => \N__33358\,
            sr => \N__49534\
        );

    \current_shift_inst.timer_s1.counter_1_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25342\,
            in1 => \N__23885\,
            in2 => \_gnd_net_\,
            in3 => \N__23866\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__49886\,
            ce => \N__33358\,
            sr => \N__49534\
        );

    \current_shift_inst.timer_s1.counter_2_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25326\,
            in1 => \N__23855\,
            in2 => \_gnd_net_\,
            in3 => \N__23839\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__49886\,
            ce => \N__33358\,
            sr => \N__49534\
        );

    \current_shift_inst.timer_s1.counter_3_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25343\,
            in1 => \N__23828\,
            in2 => \_gnd_net_\,
            in3 => \N__23812\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__49886\,
            ce => \N__33358\,
            sr => \N__49534\
        );

    \current_shift_inst.timer_s1.counter_4_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25327\,
            in1 => \N__23804\,
            in2 => \_gnd_net_\,
            in3 => \N__23785\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__49886\,
            ce => \N__33358\,
            sr => \N__49534\
        );

    \current_shift_inst.timer_s1.counter_5_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25344\,
            in1 => \N__23777\,
            in2 => \_gnd_net_\,
            in3 => \N__23758\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__49886\,
            ce => \N__33358\,
            sr => \N__49534\
        );

    \current_shift_inst.timer_s1.counter_6_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25328\,
            in1 => \N__23744\,
            in2 => \_gnd_net_\,
            in3 => \N__23728\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__49886\,
            ce => \N__33358\,
            sr => \N__49534\
        );

    \current_shift_inst.timer_s1.counter_7_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25345\,
            in1 => \N__24122\,
            in2 => \_gnd_net_\,
            in3 => \N__24106\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__49886\,
            ce => \N__33358\,
            sr => \N__49534\
        );

    \current_shift_inst.timer_s1.counter_8_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25324\,
            in1 => \N__24098\,
            in2 => \_gnd_net_\,
            in3 => \N__24079\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__49879\,
            ce => \N__33356\,
            sr => \N__49538\
        );

    \current_shift_inst.timer_s1.counter_9_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25332\,
            in1 => \N__24065\,
            in2 => \_gnd_net_\,
            in3 => \N__24046\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__49879\,
            ce => \N__33356\,
            sr => \N__49538\
        );

    \current_shift_inst.timer_s1.counter_10_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25321\,
            in1 => \N__24041\,
            in2 => \_gnd_net_\,
            in3 => \N__24025\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__49879\,
            ce => \N__33356\,
            sr => \N__49538\
        );

    \current_shift_inst.timer_s1.counter_11_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25329\,
            in1 => \N__24017\,
            in2 => \_gnd_net_\,
            in3 => \N__23998\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__49879\,
            ce => \N__33356\,
            sr => \N__49538\
        );

    \current_shift_inst.timer_s1.counter_12_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25322\,
            in1 => \N__23990\,
            in2 => \_gnd_net_\,
            in3 => \N__23971\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__49879\,
            ce => \N__33356\,
            sr => \N__49538\
        );

    \current_shift_inst.timer_s1.counter_13_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25330\,
            in1 => \N__23963\,
            in2 => \_gnd_net_\,
            in3 => \N__23944\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__49879\,
            ce => \N__33356\,
            sr => \N__49538\
        );

    \current_shift_inst.timer_s1.counter_14_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25323\,
            in1 => \N__23933\,
            in2 => \_gnd_net_\,
            in3 => \N__23917\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__49879\,
            ce => \N__33356\,
            sr => \N__49538\
        );

    \current_shift_inst.timer_s1.counter_15_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25331\,
            in1 => \N__24350\,
            in2 => \_gnd_net_\,
            in3 => \N__24334\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__49879\,
            ce => \N__33356\,
            sr => \N__49538\
        );

    \current_shift_inst.timer_s1.counter_16_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25311\,
            in1 => \N__24326\,
            in2 => \_gnd_net_\,
            in3 => \N__24307\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_23_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__49871\,
            ce => \N__33357\,
            sr => \N__49542\
        );

    \current_shift_inst.timer_s1.counter_17_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25315\,
            in1 => \N__24296\,
            in2 => \_gnd_net_\,
            in3 => \N__24277\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__49871\,
            ce => \N__33357\,
            sr => \N__49542\
        );

    \current_shift_inst.timer_s1.counter_18_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25312\,
            in1 => \N__24272\,
            in2 => \_gnd_net_\,
            in3 => \N__24256\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__49871\,
            ce => \N__33357\,
            sr => \N__49542\
        );

    \current_shift_inst.timer_s1.counter_19_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25316\,
            in1 => \N__24248\,
            in2 => \_gnd_net_\,
            in3 => \N__24229\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__49871\,
            ce => \N__33357\,
            sr => \N__49542\
        );

    \current_shift_inst.timer_s1.counter_20_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25313\,
            in1 => \N__24221\,
            in2 => \_gnd_net_\,
            in3 => \N__24202\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__49871\,
            ce => \N__33357\,
            sr => \N__49542\
        );

    \current_shift_inst.timer_s1.counter_21_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25317\,
            in1 => \N__24194\,
            in2 => \_gnd_net_\,
            in3 => \N__24175\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__49871\,
            ce => \N__33357\,
            sr => \N__49542\
        );

    \current_shift_inst.timer_s1.counter_22_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25314\,
            in1 => \N__24164\,
            in2 => \_gnd_net_\,
            in3 => \N__24148\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__49871\,
            ce => \N__33357\,
            sr => \N__49542\
        );

    \current_shift_inst.timer_s1.counter_23_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25318\,
            in1 => \N__24143\,
            in2 => \_gnd_net_\,
            in3 => \N__24127\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__49871\,
            ce => \N__33357\,
            sr => \N__49542\
        );

    \current_shift_inst.timer_s1.counter_24_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25307\,
            in1 => \N__24503\,
            in2 => \_gnd_net_\,
            in3 => \N__24484\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_24_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__49867\,
            ce => \N__33341\,
            sr => \N__49543\
        );

    \current_shift_inst.timer_s1.counter_25_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25319\,
            in1 => \N__24473\,
            in2 => \_gnd_net_\,
            in3 => \N__24454\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__49867\,
            ce => \N__33341\,
            sr => \N__49543\
        );

    \current_shift_inst.timer_s1.counter_26_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25308\,
            in1 => \N__24449\,
            in2 => \_gnd_net_\,
            in3 => \N__24433\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__49867\,
            ce => \N__33341\,
            sr => \N__49543\
        );

    \current_shift_inst.timer_s1.counter_27_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25320\,
            in1 => \N__24425\,
            in2 => \_gnd_net_\,
            in3 => \N__24406\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__49867\,
            ce => \N__33341\,
            sr => \N__49543\
        );

    \current_shift_inst.timer_s1.counter_28_LC_8_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25309\,
            in1 => \N__24399\,
            in2 => \_gnd_net_\,
            in3 => \N__24385\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__49867\,
            ce => \N__33341\,
            sr => \N__49543\
        );

    \current_shift_inst.timer_s1.counter_29_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24375\,
            in1 => \N__25310\,
            in2 => \_gnd_net_\,
            in3 => \N__24382\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49867\,
            ce => \N__33341\,
            sr => \N__49543\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29338\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__29262\,
            in1 => \N__29416\,
            in2 => \_gnd_net_\,
            in3 => \N__24570\,
            lcout => \current_shift_inst.PI_CTRL.un1_enablelt3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24553\,
            in1 => \N__24613\,
            in2 => \N__24520\,
            in3 => \N__24541\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38036\,
            in1 => \N__29203\,
            in2 => \N__38178\,
            in3 => \N__29998\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110101"
        )
    port map (
            in0 => \N__29566\,
            in1 => \N__24547\,
            in2 => \N__24532\,
            in3 => \N__34797\,
            lcout => \current_shift_inst.PI_CTRL.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33950\,
            in2 => \_gnd_net_\,
            in3 => \N__29633\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__38095\,
            in1 => \N__37100\,
            in2 => \N__24535\,
            in3 => \N__29328\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27175\,
            in2 => \_gnd_net_\,
            in3 => \N__33863\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24601\,
            in1 => \N__24619\,
            in2 => \N__24523\,
            in3 => \N__24595\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29784\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35446\,
            in1 => \N__35634\,
            in2 => \N__29842\,
            in3 => \N__35104\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34085\,
            in1 => \N__29785\,
            in2 => \N__25379\,
            in3 => \N__37444\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33703\,
            in1 => \N__35265\,
            in2 => \N__29482\,
            in3 => \N__34006\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27133\,
            in1 => \N__30304\,
            in2 => \N__33812\,
            in3 => \N__29703\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34060\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33702\,
            in1 => \N__35266\,
            in2 => \N__29483\,
            in3 => \N__34007\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35103\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25375\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33949\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__37439\,
            in1 => \N__37283\,
            in2 => \N__37665\,
            in3 => \N__27046\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49461\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__37282\,
            in1 => \N__37440\,
            in2 => \N__27034\,
            in3 => \N__37602\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49461\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30058\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49944\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33753\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49944\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30034\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49944\,
            ce => 'H',
            sr => \N__49468\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35018\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49944\,
            ce => 'H',
            sr => \N__49468\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24631\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32853\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32642\,
            in1 => \N__32090\,
            in2 => \N__24724\,
            in3 => \N__24683\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000101"
        )
    port map (
            in0 => \N__24763\,
            in1 => \N__24782\,
            in2 => \N__32139\,
            in3 => \N__32645\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__32644\,
            in1 => \N__32092\,
            in2 => \N__24786\,
            in3 => \N__24762\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__32088\,
            in1 => \N__32640\,
            in2 => \N__27352\,
            in3 => \N__27299\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32641\,
            in1 => \N__32089\,
            in2 => \N__30765\,
            in3 => \N__30713\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__32086\,
            in1 => \N__27432\,
            in2 => \N__24838\,
            in3 => \N__24817\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32639\,
            in1 => \N__32087\,
            in2 => \N__30850\,
            in3 => \N__30791\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__32091\,
            in1 => \N__24723\,
            in2 => \N__24688\,
            in3 => \N__32643\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32717\,
            in1 => \N__31990\,
            in2 => \N__30535\,
            in3 => \N__30485\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__31992\,
            in1 => \N__32719\,
            in2 => \N__30939\,
            in3 => \N__30884\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__30657\,
            in1 => \N__24833\,
            in2 => \_gnd_net_\,
            in3 => \N__24812\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__31987\,
            in1 => \N__32721\,
            in2 => \N__25879\,
            in3 => \N__25923\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32720\,
            in1 => \N__31993\,
            in2 => \N__31369\,
            in3 => \N__31301\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__31988\,
            in1 => \N__30963\,
            in2 => \N__31014\,
            in3 => \N__32722\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__32716\,
            in1 => \N__31442\,
            in2 => \N__31423\,
            in3 => \N__31989\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__31991\,
            in1 => \N__32718\,
            in2 => \N__26137\,
            in3 => \N__26094\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__32114\,
            in1 => \N__32637\,
            in2 => \N__25971\,
            in3 => \N__25994\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__26133\,
            in1 => \N__30624\,
            in2 => \_gnd_net_\,
            in3 => \N__26093\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__32117\,
            in1 => \N__32634\,
            in2 => \N__31243\,
            in3 => \N__31262\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32635\,
            in1 => \N__32118\,
            in2 => \N__31564\,
            in3 => \N__31508\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__32119\,
            in1 => \N__31652\,
            in2 => \N__31612\,
            in3 => \N__32636\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32638\,
            in1 => \N__32115\,
            in2 => \N__26077\,
            in3 => \N__26021\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30623\,
            in1 => \N__31001\,
            in2 => \_gnd_net_\,
            in3 => \N__30962\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32633\,
            in1 => \N__32116\,
            in2 => \N__24904\,
            in3 => \N__24858\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__32122\,
            in1 => \N__24954\,
            in2 => \N__24925\,
            in3 => \N__32673\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__24955\,
            in1 => \N__24921\,
            in2 => \N__32715\,
            in3 => \N__32123\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32120\,
            in1 => \N__24953\,
            in2 => \_gnd_net_\,
            in3 => \N__24915\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__32672\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32124\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__32121\,
            in1 => \N__32677\,
            in2 => \N__24859\,
            in3 => \N__24900\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30630\,
            in1 => \N__24899\,
            in2 => \_gnd_net_\,
            in3 => \N__24854\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27666\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49909\,
            ce => \N__27633\,
            sr => \N__49510\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27995\,
            in2 => \N__26541\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28070\,
            in2 => \N__25012\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25000\,
            in2 => \N__28164\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28074\,
            in2 => \N__24994\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24985\,
            in2 => \N__28165\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28078\,
            in2 => \N__24979\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24970\,
            in2 => \N__28166\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28082\,
            in2 => \N__24964\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28179\,
            in2 => \N__25066\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25057\,
            in2 => \N__28269\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28167\,
            in2 => \N__25048\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30463\,
            in2 => \N__28266\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28171\,
            in2 => \N__25036\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25024\,
            in2 => \N__28267\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28175\,
            in2 => \N__26389\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25018\,
            in2 => \N__28268\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28183\,
            in2 => \N__25120\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25111\,
            in2 => \N__28270\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28187\,
            in2 => \N__25105\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25096\,
            in2 => \N__28271\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28191\,
            in2 => \N__26398\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25090\,
            in2 => \N__28272\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28195\,
            in2 => \N__25081\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25072\,
            in2 => \N__28273\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28199\,
            in2 => \N__25204\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25195\,
            in2 => \N__28274\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28203\,
            in2 => \N__25189\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25180\,
            in2 => \N__28275\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28207\,
            in2 => \N__25171\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25156\,
            in2 => \N__28276\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28211\,
            in2 => \N__25150\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32147\,
            in2 => \_gnd_net_\,
            in3 => \N__25135\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41261\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49880\,
            ce => 'H',
            sr => \N__49530\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34879\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35884\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49851\,
            ce => 'H',
            sr => \N__49544\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__37673\,
            in1 => \N__37307\,
            in2 => \_gnd_net_\,
            in3 => \N__26707\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49963\,
            ce => 'H',
            sr => \N__49414\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25210\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49959\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29420\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29193\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29481\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29261\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29559\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110011111110"
        )
    port map (
            in0 => \N__37230\,
            in1 => \N__37456\,
            in2 => \N__37706\,
            in3 => \N__26647\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49430\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110101110"
        )
    port map (
            in0 => \N__37453\,
            in1 => \N__37231\,
            in2 => \N__26743\,
            in3 => \N__37686\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49430\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110101110"
        )
    port map (
            in0 => \N__37454\,
            in1 => \N__37232\,
            in2 => \N__26926\,
            in3 => \N__37687\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49430\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110101110"
        )
    port map (
            in0 => \N__37455\,
            in1 => \N__37233\,
            in2 => \N__26857\,
            in3 => \N__37688\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49949\,
            ce => 'H',
            sr => \N__49430\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__37269\,
            in1 => \N__37452\,
            in2 => \N__26947\,
            in3 => \N__37629\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => 'H',
            sr => \N__49437\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__37447\,
            in1 => \N__37272\,
            in2 => \N__37671\,
            in3 => \N__26980\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => 'H',
            sr => \N__49437\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__37267\,
            in1 => \N__37450\,
            in2 => \N__26869\,
            in3 => \N__37628\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => 'H',
            sr => \N__49437\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__37445\,
            in1 => \N__37270\,
            in2 => \N__37669\,
            in3 => \N__26761\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => 'H',
            sr => \N__49437\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__37266\,
            in1 => \N__37449\,
            in2 => \N__26905\,
            in3 => \N__37627\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => 'H',
            sr => \N__49437\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__37448\,
            in1 => \N__37273\,
            in2 => \N__37672\,
            in3 => \N__26971\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => 'H',
            sr => \N__49437\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__37268\,
            in1 => \N__37451\,
            in2 => \N__26827\,
            in3 => \N__37630\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => 'H',
            sr => \N__49437\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__37446\,
            in1 => \N__37271\,
            in2 => \N__37670\,
            in3 => \N__26890\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => 'H',
            sr => \N__49437\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33258\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49448\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111101010100"
        )
    port map (
            in0 => \N__26989\,
            in1 => \N__37308\,
            in2 => \N__37708\,
            in3 => \N__37442\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49448\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49448\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010111"
        )
    port map (
            in0 => \N__26806\,
            in1 => \N__37693\,
            in2 => \N__37325\,
            in3 => \N__37443\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49448\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33288\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49448\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011101010100"
        )
    port map (
            in0 => \N__27016\,
            in1 => \N__37692\,
            in2 => \N__37324\,
            in3 => \N__37441\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => 'H',
            sr => \N__49448\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49456\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__37315\,
            in1 => \N__37438\,
            in2 => \N__27202\,
            in3 => \N__37682\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49456\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37932\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49456\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30090\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49456\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__28998\,
            in1 => \N__35366\,
            in2 => \_gnd_net_\,
            in3 => \N__29059\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49919\,
            ce => 'H',
            sr => \N__49469\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__32881\,
            in1 => \N__26223\,
            in2 => \_gnd_net_\,
            in3 => \N__26185\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49919\,
            ce => 'H',
            sr => \N__49469\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27925\,
            in2 => \N__27942\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27422\,
            in2 => \N__25447\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32598\,
            in2 => \N__27541\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25438\,
            in2 => \N__32669\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32602\,
            in2 => \N__25432\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25624\,
            in2 => \N__32670\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32606\,
            in2 => \N__25618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25609\,
            in2 => \N__32671\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32330\,
            in2 => \N__25603\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25594\,
            in2 => \N__32525\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32334\,
            in2 => \N__25588\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25579\,
            in2 => \N__32526\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32338\,
            in2 => \N__25573\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25564\,
            in2 => \N__32527\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32342\,
            in2 => \N__25660\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25651\,
            in2 => \N__32528\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32362\,
            in2 => \N__26236\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31024\,
            in2 => \N__32533\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32366\,
            in2 => \N__25645\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30859\,
            in2 => \N__32534\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32370\,
            in2 => \N__31111\,
            in3 => \N__25636\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25633\,
            in2 => \N__32535\,
            in3 => \N__25627\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32374\,
            in2 => \N__25771\,
            in3 => \N__25759\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25756\,
            in2 => \N__32536\,
            in3 => \N__25750\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32431\,
            in2 => \N__25747\,
            in3 => \N__25738\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25735\,
            in2 => \N__32585\,
            in3 => \N__25726\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32435\,
            in2 => \N__25723\,
            in3 => \N__25711\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27214\,
            in2 => \N__32586\,
            in3 => \N__25708\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32439\,
            in2 => \N__25705\,
            in3 => \N__25693\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25690\,
            in2 => \N__32587\,
            in3 => \N__25681\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32443\,
            in2 => \N__25678\,
            in3 => \N__25663\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__32444\,
            in1 => \N__32128\,
            in2 => \_gnd_net_\,
            in3 => \N__26140\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32015\,
            in1 => \N__26132\,
            in2 => \N__32653\,
            in3 => \N__26101\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__31063\,
            in1 => \N__32018\,
            in2 => \N__31099\,
            in3 => \N__32571\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__26310\,
            in1 => \N__32017\,
            in2 => \N__26272\,
            in3 => \N__32570\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__32572\,
            in1 => \N__26076\,
            in2 => \N__32107\,
            in3 => \N__26032\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__25999\,
            in1 => \N__32569\,
            in2 => \N__25975\,
            in3 => \N__32016\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32014\,
            in1 => \N__25924\,
            in2 => \N__32654\,
            in3 => \N__25875\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31232\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__25831\,
            in1 => \N__32111\,
            in2 => \N__32724\,
            in3 => \N__25798\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32693\,
            in1 => \N__32112\,
            in2 => \N__26488\,
            in3 => \N__26446\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__32113\,
            in1 => \N__32701\,
            in2 => \N__27996\,
            in3 => \N__26419\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__31182\,
            in1 => \N__30653\,
            in2 => \_gnd_net_\,
            in3 => \N__31137\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30652\,
            in1 => \N__31352\,
            in2 => \_gnd_net_\,
            in3 => \N__31311\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__26377\,
            in1 => \N__32110\,
            in2 => \N__32723\,
            in3 => \N__26341\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__32109\,
            in1 => \N__32700\,
            in2 => \N__26314\,
            in3 => \N__26265\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__32892\,
            in1 => \N__26224\,
            in2 => \_gnd_net_\,
            in3 => \N__26181\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_398_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36228\,
            in2 => \_gnd_net_\,
            in3 => \N__36181\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32891\,
            in2 => \_gnd_net_\,
            in3 => \N__26180\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_397_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__26542\,
            in1 => \N__28212\,
            in2 => \_gnd_net_\,
            in3 => \N__26512\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27659\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49868\,
            ce => \N__27626\,
            sr => \N__49524\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28927\,
            in2 => \N__28720\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43124\,
            in1 => \N__27891\,
            in2 => \_gnd_net_\,
            in3 => \N__26506\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49526\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__43121\,
            in1 => \N__28578\,
            in2 => \N__28744\,
            in3 => \N__26503\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49526\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43125\,
            in1 => \N__28554\,
            in2 => \_gnd_net_\,
            in3 => \N__26500\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49526\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43122\,
            in1 => \N__28533\,
            in2 => \_gnd_net_\,
            in3 => \N__26497\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49526\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43126\,
            in1 => \N__28506\,
            in2 => \_gnd_net_\,
            in3 => \N__26494\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49526\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43123\,
            in1 => \N__28482\,
            in2 => \_gnd_net_\,
            in3 => \N__26491\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49526\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43127\,
            in1 => \N__28461\,
            in2 => \_gnd_net_\,
            in3 => \N__26569\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49526\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43096\,
            in1 => \N__28434\,
            in2 => \_gnd_net_\,
            in3 => \N__26566\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49858\,
            ce => 'H',
            sr => \N__49531\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43089\,
            in1 => \N__28410\,
            in2 => \_gnd_net_\,
            in3 => \N__26563\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49858\,
            ce => 'H',
            sr => \N__49531\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43093\,
            in1 => \N__28695\,
            in2 => \_gnd_net_\,
            in3 => \N__26560\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49858\,
            ce => 'H',
            sr => \N__49531\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43090\,
            in1 => \N__28671\,
            in2 => \_gnd_net_\,
            in3 => \N__26557\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49858\,
            ce => 'H',
            sr => \N__49531\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43094\,
            in1 => \N__28647\,
            in2 => \_gnd_net_\,
            in3 => \N__26554\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49858\,
            ce => 'H',
            sr => \N__49531\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43091\,
            in1 => \N__28623\,
            in2 => \_gnd_net_\,
            in3 => \N__26551\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49858\,
            ce => 'H',
            sr => \N__49531\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43095\,
            in1 => \N__28599\,
            in2 => \_gnd_net_\,
            in3 => \N__26548\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49858\,
            ce => 'H',
            sr => \N__49531\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43092\,
            in1 => \N__42708\,
            in2 => \_gnd_net_\,
            in3 => \N__26545\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49858\,
            ce => 'H',
            sr => \N__49531\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43139\,
            in1 => \N__42675\,
            in2 => \_gnd_net_\,
            in3 => \N__26596\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49535\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43132\,
            in1 => \N__42842\,
            in2 => \_gnd_net_\,
            in3 => \N__26593\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49535\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43140\,
            in1 => \N__42870\,
            in2 => \_gnd_net_\,
            in3 => \N__26590\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49535\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43133\,
            in1 => \N__28870\,
            in2 => \_gnd_net_\,
            in3 => \N__26587\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49535\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43141\,
            in1 => \N__28882\,
            in2 => \_gnd_net_\,
            in3 => \N__26584\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49535\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43134\,
            in1 => \N__28837\,
            in2 => \_gnd_net_\,
            in3 => \N__26581\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49535\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43142\,
            in1 => \N__28849\,
            in2 => \_gnd_net_\,
            in3 => \N__26578\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49535\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43135\,
            in1 => \N__28804\,
            in2 => \_gnd_net_\,
            in3 => \N__26575\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49535\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43128\,
            in1 => \N__28816\,
            in2 => \_gnd_net_\,
            in3 => \N__26572\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_10_25_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49852\,
            ce => 'H',
            sr => \N__49539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43136\,
            in1 => \N__28771\,
            in2 => \_gnd_net_\,
            in3 => \N__26614\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49852\,
            ce => 'H',
            sr => \N__49539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43129\,
            in1 => \N__28783\,
            in2 => \_gnd_net_\,
            in3 => \N__26611\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49852\,
            ce => 'H',
            sr => \N__49539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43137\,
            in1 => \N__29143\,
            in2 => \_gnd_net_\,
            in3 => \N__26608\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49852\,
            ce => 'H',
            sr => \N__49539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43130\,
            in1 => \N__29155\,
            in2 => \_gnd_net_\,
            in3 => \N__26605\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49852\,
            ce => 'H',
            sr => \N__49539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43138\,
            in1 => \N__29088\,
            in2 => \_gnd_net_\,
            in3 => \N__26602\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49852\,
            ce => 'H',
            sr => \N__49539\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43131\,
            in1 => \N__29114\,
            in2 => \_gnd_net_\,
            in3 => \N__26599\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49852\,
            ce => 'H',
            sr => \N__49539\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34774\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__37983\,
            in1 => \N__34775\,
            in2 => \N__33463\,
            in3 => \N__30121\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29614\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101100011011"
        )
    port map (
            in0 => \N__37707\,
            in1 => \N__37499\,
            in2 => \N__26629\,
            in3 => \N__37303\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49953\,
            ce => 'H',
            sr => \N__49415\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37091\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29652\,
            in2 => \N__29656\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29373\,
            in2 => \N__29356\,
            in3 => \N__26719\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26716\,
            in2 => \N__29389\,
            in3 => \N__26698\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26695\,
            in2 => \N__29224\,
            in3 => \N__26680\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26677\,
            in2 => \N__26668\,
            in3 => \N__26656\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26653\,
            in2 => \N__29533\,
            in3 => \N__26641\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29593\,
            in2 => \N__26638\,
            in3 => \N__26617\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26818\,
            in2 => \N__29290\,
            in3 => \N__26797\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26794\,
            in2 => \N__29164\,
            in3 => \N__26782\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26779\,
            in2 => \N__35146\,
            in3 => \N__26770\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35599\,
            in2 => \N__29281\,
            in3 => \N__26767\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29503\,
            in2 => \N__29524\,
            in3 => \N__26764\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27103\,
            in2 => \N__35230\,
            in3 => \N__26755\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26752\,
            in2 => \N__29755\,
            in3 => \N__26734\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29497\,
            in2 => \N__29512\,
            in3 => \N__26731\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26932\,
            in2 => \N__29173\,
            in3 => \N__26917\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26914\,
            in2 => \N__29443\,
            in3 => \N__26896\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35317\,
            in2 => \N__37729\,
            in3 => \N__26893\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33676\,
            in2 => \N__29665\,
            in3 => \N__26884\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26881\,
            in2 => \N__35056\,
            in3 => \N__26860\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35608\,
            in2 => \N__29746\,
            in3 => \N__26848\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29938\,
            in2 => \N__29947\,
            in3 => \N__26845\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29725\,
            in2 => \N__33769\,
            in3 => \N__26842\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29803\,
            in2 => \N__26839\,
            in3 => \N__27049\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27394\,
            in2 => \N__29956\,
            in3 => \N__27037\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34120\,
            in2 => \N__35398\,
            in3 => \N__27022\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27079\,
            in2 => \N__29737\,
            in3 => \N__27019\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27073\,
            in2 => \N__29677\,
            in3 => \N__27007\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34039\,
            in2 => \N__27004\,
            in3 => \N__26983\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27092\,
            in2 => \N__27112\,
            in3 => \N__26974\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27094\,
            in2 => \N__27157\,
            in3 => \N__26965\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27093\,
            in2 => \N__26962\,
            in3 => \N__26935\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un13_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un13_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37460\,
            in1 => \N__37838\,
            in2 => \_gnd_net_\,
            in3 => \N__27205\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27189\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27140\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35273\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37837\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30291\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29704\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27064\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49920\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__35365\,
            in1 => \N__29055\,
            in2 => \_gnd_net_\,
            in3 => \N__28997\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_400_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29999\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__27385\,
            in1 => \N__27856\,
            in2 => \_gnd_net_\,
            in3 => \N__32850\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27376\,
            in3 => \N__30257\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => 'H',
            sr => \N__49462\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32851\,
            lcout => \current_shift_inst.N_1474_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__32852\,
            in1 => \N__27373\,
            in2 => \_gnd_net_\,
            in3 => \N__27829\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__28351\,
            in1 => \N__27364\,
            in2 => \_gnd_net_\,
            in3 => \N__32848\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__31957\,
            in1 => \N__27348\,
            in2 => \N__32668\,
            in3 => \N__27304\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__27280\,
            in1 => \N__32445\,
            in2 => \N__27238\,
            in3 => \N__31956\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000101"
        )
    port map (
            in0 => \N__27279\,
            in1 => \N__27234\,
            in2 => \N__32025\,
            in3 => \N__32446\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27670\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49905\,
            ce => \N__27632\,
            sr => \N__49478\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__31952\,
            in1 => \N__32447\,
            in2 => \N__27574\,
            in3 => \N__27601\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__27600\,
            in1 => \N__27570\,
            in2 => \N__32588\,
            in3 => \N__31950\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__31951\,
            in1 => \N__27502\,
            in2 => \_gnd_net_\,
            in3 => \N__27493\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27532\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__31949\,
            in1 => \_gnd_net_\,
            in2 => \N__27496\,
            in3 => \N__27492\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27924\,
            in2 => \N__27460\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27991\,
            in1 => \N__27418\,
            in2 => \N__27451\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32318\,
            in2 => \N__27727\,
            in3 => \N__27990\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30772\,
            in2 => \N__32522\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32322\,
            in2 => \N__27718\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30691\,
            in2 => \N__32523\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32326\,
            in2 => \N__27706\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27691\,
            in2 => \N__32524\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32346\,
            in2 => \N__27679\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30946\,
            in2 => \N__32529\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32350\,
            in2 => \N__31378\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27775\,
            in2 => \N__32530\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32354\,
            in2 => \N__27766\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30865\,
            in2 => \N__32531\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32358\,
            in2 => \N__31282\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27757\,
            in2 => \N__32532\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32537\,
            in2 => \N__27751\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27742\,
            in2 => \N__32646\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32541\,
            in2 => \N__27736\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31759\,
            in2 => \N__32647\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32545\,
            in2 => \N__27871\,
            in3 => \N__27844\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27841\,
            in2 => \N__32648\,
            in3 => \N__27820\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32549\,
            in2 => \N__31198\,
            in3 => \N__27817\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31489\,
            in2 => \N__32649\,
            in3 => \N__27814\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32553\,
            in2 => \N__31576\,
            in3 => \N__27811\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27808\,
            in2 => \N__32650\,
            in3 => \N__27802\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32557\,
            in2 => \N__27799\,
            in3 => \N__27790\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27787\,
            in2 => \N__32651\,
            in3 => \N__27778\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32561\,
            in2 => \N__28387\,
            in3 => \N__28372\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28369\,
            in2 => \N__32652\,
            in3 => \N__28363\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32565\,
            in2 => \N__28360\,
            in3 => \N__28342\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__28339\,
            in1 => \N__28327\,
            in2 => \N__32849\,
            in3 => \N__28318\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__47112\,
            in1 => \N__34518\,
            in2 => \_gnd_net_\,
            in3 => \N__42213\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49873\,
            ce => \N__49120\,
            sr => \N__49511\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__28220\,
            in1 => \N__27972\,
            in2 => \_gnd_net_\,
            in3 => \N__27943\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33166\,
            in2 => \N__27904\,
            in3 => \N__28719\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27877\,
            in2 => \N__31726\,
            in3 => \N__27895\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31747\,
            in2 => \N__28564\,
            in3 => \N__28579\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28540\,
            in2 => \N__31714\,
            in3 => \N__28555\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31702\,
            in2 => \N__28519\,
            in3 => \N__28534\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31735\,
            in2 => \N__28492\,
            in3 => \N__28507\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28483\,
            in1 => \N__28468\,
            in2 => \N__33175\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28462\,
            in1 => \N__32734\,
            in2 => \N__28447\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43165\,
            in2 => \N__28420\,
            in3 => \N__28438\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43276\,
            in2 => \N__28396\,
            in3 => \N__28411\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43234\,
            in2 => \N__28681\,
            in3 => \N__28696\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43195\,
            in2 => \N__28657\,
            in3 => \N__28672\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43180\,
            in2 => \N__28633\,
            in3 => \N__28648\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28624\,
            in1 => \N__43324\,
            in2 => \N__28609\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28600\,
            in1 => \N__28585\,
            in2 => \N__34684\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42661\,
            in2 => \N__42739\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28891\,
            in2 => \N__42820\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28858\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28825\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28792\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28759\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29131\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29068\,
            in2 => \N__29122\,
            in3 => \N__28750\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28747\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010011101110"
        )
    port map (
            in0 => \N__28920\,
            in1 => \N__28732\,
            in2 => \N__28906\,
            in3 => \N__33086\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \N__49527\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28919\,
            in2 => \_gnd_net_\,
            in3 => \N__28938\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__33061\,
            in1 => \N__33084\,
            in2 => \_gnd_net_\,
            in3 => \N__28731\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__43042\,
            in1 => \N__28939\,
            in2 => \N__28723\,
            in3 => \N__28718\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \N__49527\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111111"
        )
    port map (
            in0 => \N__29089\,
            in1 => \N__29115\,
            in2 => \N__28951\,
            in3 => \N__33085\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28930\,
            in3 => \N__28918\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110100001000"
        )
    port map (
            in0 => \N__28921\,
            in1 => \N__33087\,
            in2 => \N__28905\,
            in3 => \N__44624\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \N__49527\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__43345\,
            in1 => \N__42866\,
            in2 => \N__42846\,
            in3 => \N__42898\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28881\,
            in2 => \_gnd_net_\,
            in3 => \N__28869\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__28848\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28836\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28815\,
            in2 => \_gnd_net_\,
            in3 => \N__28803\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28782\,
            in2 => \_gnd_net_\,
            in3 => \N__28770\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29154\,
            in2 => \_gnd_net_\,
            in3 => \N__29142\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_df28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29113\,
            in2 => \_gnd_net_\,
            in3 => \N__29087\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29048\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29020\,
            ce => 'H',
            sr => \N__49536\
        );

    \delay_measurement_inst.start_timer_tr_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29047\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29019\,
            ce => 'H',
            sr => \N__49540\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35383\,
            in2 => \_gnd_net_\,
            in3 => \N__29008\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_399_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30120\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30146\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29912\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29882\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__37878\,
            in1 => \N__29430\,
            in2 => \N__29887\,
            in3 => \N__33184\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__29377\,
            in1 => \N__37877\,
            in2 => \N__29917\,
            in3 => \N__33199\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__37882\,
            in1 => \N__29339\,
            in2 => \N__33415\,
            in3 => \N__30057\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__38096\,
            in1 => \N__37883\,
            in2 => \N__33754\,
            in3 => \N__33376\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \N__29266\,
            in1 => \N__30147\,
            in2 => \N__37942\,
            in3 => \N__33478\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30086\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30056\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__33546\,
            in1 => \N__29214\,
            in2 => \N__33529\,
            in3 => \N__37974\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__37972\,
            in1 => \N__33951\,
            in2 => \N__33394\,
            in3 => \N__30033\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37969\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__37971\,
            in1 => \N__29623\,
            in2 => \N__33433\,
            in3 => \N__35020\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__29583\,
            in1 => \N__37970\,
            in2 => \N__30091\,
            in3 => \N__33442\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30032\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__35041\,
            in1 => \N__33867\,
            in2 => \N__33583\,
            in3 => \N__37973\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110101111101"
        )
    port map (
            in0 => \N__37871\,
            in1 => \N__33556\,
            in2 => \N__35494\,
            in3 => \N__38155\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33840\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38154\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__34987\,
            in1 => \N__29491\,
            in2 => \N__33514\,
            in3 => \N__37872\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__29856\,
            in1 => \N__35515\,
            in2 => \N__37941\,
            in3 => \N__33622\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__33547\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37867\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__29789\,
            in1 => \N__34144\,
            in2 => \N__37940\,
            in3 => \N__33565\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111111"
        )
    port map (
            in0 => \N__35215\,
            in1 => \N__35650\,
            in2 => \N__33664\,
            in3 => \N__37873\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__30311\,
            in1 => \N__34177\,
            in2 => \N__37944\,
            in3 => \N__33601\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33643\,
            in2 => \_gnd_net_\,
            in3 => \N__37884\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110101111101"
        )
    port map (
            in0 => \N__37888\,
            in1 => \N__33631\,
            in2 => \N__29728\,
            in3 => \N__33802\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__29719\,
            in1 => \N__37892\,
            in2 => \N__35587\,
            in3 => \N__33592\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__33716\,
            in1 => \N__35341\,
            in2 => \N__37943\,
            in3 => \N__33499\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__34109\,
            in1 => \N__30004\,
            in2 => \N__37945\,
            in3 => \N__33613\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__35308\,
            in1 => \N__37893\,
            in2 => \N__34011\,
            in3 => \N__33652\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34002\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29932\,
            in2 => \_gnd_net_\,
            in3 => \N__30235\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30220\,
            in2 => \_gnd_net_\,
            in3 => \N__29926\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30208\,
            in2 => \_gnd_net_\,
            in3 => \N__29923\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30196\,
            in2 => \_gnd_net_\,
            in3 => \N__29920\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30184\,
            in2 => \_gnd_net_\,
            in3 => \N__29890\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30172\,
            in2 => \_gnd_net_\,
            in3 => \N__29860\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30160\,
            in2 => \_gnd_net_\,
            in3 => \N__30124\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30451\,
            in2 => \_gnd_net_\,
            in3 => \N__30094\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30439\,
            in2 => \_gnd_net_\,
            in3 => \N__30064\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30427\,
            in2 => \_gnd_net_\,
            in3 => \N__30061\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30409\,
            in2 => \_gnd_net_\,
            in3 => \N__30037\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30385\,
            in2 => \_gnd_net_\,
            in3 => \N__30013\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30364\,
            in2 => \_gnd_net_\,
            in3 => \N__30010\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30337\,
            in2 => \_gnd_net_\,
            in3 => \N__30007\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30349\,
            in2 => \_gnd_net_\,
            in3 => \N__30328\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100101110"
        )
    port map (
            in0 => \N__37475\,
            in1 => \N__37681\,
            in2 => \N__30325\,
            in3 => \N__37316\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30268\,
            in2 => \N__30261\,
            in3 => \N__30262\,
            lcout => \current_shift_inst.control_input_18\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30226\,
            in2 => \_gnd_net_\,
            in3 => \N__30211\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31672\,
            in2 => \_gnd_net_\,
            in3 => \N__30199\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33022\,
            in2 => \_gnd_net_\,
            in3 => \N__30187\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32992\,
            in2 => \_gnd_net_\,
            in3 => \N__30175\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32962\,
            in2 => \_gnd_net_\,
            in3 => \N__30163\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32935\,
            in2 => \_gnd_net_\,
            in3 => \N__30151\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32905\,
            in2 => \_gnd_net_\,
            in3 => \N__30442\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32749\,
            in2 => \_gnd_net_\,
            in3 => \N__30430\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31465\,
            in2 => \_gnd_net_\,
            in3 => \N__30418\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30415\,
            in2 => \_gnd_net_\,
            in3 => \N__30400\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30397\,
            in2 => \_gnd_net_\,
            in3 => \N__30376\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30373\,
            in2 => \_gnd_net_\,
            in3 => \N__30355\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32857\,
            in2 => \_gnd_net_\,
            in3 => \N__30352\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => \current_shift_inst.control_input_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30340\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__30669\,
            in1 => \N__35844\,
            in2 => \N__30685\,
            in3 => \N__35873\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49463\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30668\,
            in2 => \_gnd_net_\,
            in3 => \N__30681\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010011110000"
        )
    port map (
            in0 => \N__35794\,
            in1 => \N__36229\,
            in2 => \N__30673\,
            in3 => \N__36141\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49463\
        );

    \phase_controller_inst2.state_1_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__35845\,
            in1 => \N__35872\,
            in2 => \_gnd_net_\,
            in3 => \N__41278\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49463\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__36140\,
            in1 => \N__36106\,
            in2 => \N__36078\,
            in3 => \N__36739\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49463\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__35740\,
            in1 => \N__38793\,
            in2 => \N__38860\,
            in3 => \N__40696\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49899\,
            ce => \N__50321\,
            sr => \N__49470\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__38792\,
            in1 => \N__41803\,
            in2 => \_gnd_net_\,
            in3 => \N__35719\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49899\,
            ce => \N__50321\,
            sr => \N__49470\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__41804\,
            in1 => \N__35683\,
            in2 => \_gnd_net_\,
            in3 => \N__38794\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49899\,
            ce => \N__50321\,
            sr => \N__49470\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__30658\,
            in1 => \N__30531\,
            in2 => \_gnd_net_\,
            in3 => \N__30486\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32451\,
            in1 => \N__31964\,
            in2 => \N__31189\,
            in3 => \N__31138\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__32453\,
            in1 => \N__31961\,
            in2 => \N__31095\,
            in3 => \N__31058\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__31960\,
            in1 => \N__32457\,
            in2 => \N__31015\,
            in3 => \N__30970\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32452\,
            in1 => \N__31962\,
            in2 => \N__30940\,
            in3 => \N__30892\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__31963\,
            in1 => \N__32454\,
            in2 => \N__31804\,
            in3 => \N__31830\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32455\,
            in1 => \N__31958\,
            in2 => \N__30849\,
            in3 => \N__30799\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__31959\,
            in1 => \N__32456\,
            in2 => \N__30766\,
            in3 => \N__30718\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36180\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49887\,
            ce => 'H',
            sr => \N__49485\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110000001100"
        )
    port map (
            in0 => \N__50058\,
            in1 => \N__34649\,
            in2 => \N__50037\,
            in3 => \N__50107\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49887\,
            ce => 'H',
            sr => \N__49485\
        );

    \phase_controller_inst1.state_4_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__33140\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44532\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49887\,
            ce => 'H',
            sr => \N__49485\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__32137\,
            in1 => \N__31657\,
            in2 => \N__31608\,
            in3 => \N__32594\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__32593\,
            in1 => \N__32136\,
            in2 => \N__31563\,
            in3 => \N__31516\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__31483\,
            in1 => \N__31477\,
            in2 => \_gnd_net_\,
            in3 => \N__32828\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__32595\,
            in1 => \N__32132\,
            in2 => \N__31456\,
            in3 => \N__31419\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__32133\,
            in1 => \N__32596\,
            in2 => \N__31368\,
            in3 => \N__31312\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__32592\,
            in1 => \N__32135\,
            in2 => \N__31273\,
            in3 => \N__31239\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39516\,
            in1 => \N__42547\,
            in2 => \N__39493\,
            in3 => \N__42525\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__32597\,
            in1 => \N__32134\,
            in2 => \N__31837\,
            in3 => \N__31803\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111010"
        )
    port map (
            in0 => \N__46015\,
            in1 => \N__39241\,
            in2 => \N__34609\,
            in3 => \N__45547\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31753\,
            in3 => \N__45370\,
            lcout => \elapsed_time_ns_1_RNIRB3CP1_0_3\,
            ltout => \elapsed_time_ns_1_RNIRB3CP1_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__42280\,
            in1 => \N__42201\,
            in2 => \N__31750\,
            in3 => \N__34483\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => \N__43150\,
            sr => \N__49500\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__47088\,
            in1 => \N__45964\,
            in2 => \N__42215\,
            in3 => \N__42283\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => \N__43150\,
            sr => \N__49500\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__42279\,
            in1 => \N__47085\,
            in2 => \N__34702\,
            in3 => \N__42200\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => \N__43150\,
            sr => \N__49500\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__47086\,
            in1 => \N__42282\,
            in2 => \N__42214\,
            in3 => \N__39303\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => \N__43150\,
            sr => \N__49500\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__42281\,
            in1 => \N__47087\,
            in2 => \N__42313\,
            in3 => \N__42202\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49872\,
            ce => \N__43150\,
            sr => \N__49500\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31693\,
            in1 => \N__31681\,
            in2 => \_gnd_net_\,
            in3 => \N__32821\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__32823\,
            in1 => \N__33043\,
            in2 => \_gnd_net_\,
            in3 => \N__33031\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__33010\,
            in1 => \N__32998\,
            in2 => \_gnd_net_\,
            in3 => \N__32824\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100100111"
        )
    port map (
            in0 => \N__32826\,
            in1 => \N__32983\,
            in2 => \N__32977\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__32953\,
            in1 => \N__32947\,
            in2 => \_gnd_net_\,
            in3 => \N__32822\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__32825\,
            in1 => \N__32923\,
            in2 => \_gnd_net_\,
            in3 => \N__32917\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32893\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__32827\,
            in1 => \N__32767\,
            in2 => \_gnd_net_\,
            in3 => \N__32755\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__47098\,
            in1 => \N__42204\,
            in2 => \_gnd_net_\,
            in3 => \N__34519\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => \N__43144\,
            sr => \N__49512\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__47097\,
            in1 => \N__42203\,
            in2 => \N__38323\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => \N__43144\,
            sr => \N__49512\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__34534\,
            in1 => \N__42284\,
            in2 => \N__34720\,
            in3 => \N__34735\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49862\,
            ce => \N__43144\,
            sr => \N__49512\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38246\,
            in2 => \_gnd_net_\,
            in3 => \N__38295\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a2_1_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33149\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44541\,
            lcout => state_ns_i_a2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33066\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \N__49522\
        );

    \phase_controller_inst1.state_1_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__33367\,
            in1 => \N__44601\,
            in2 => \_gnd_net_\,
            in3 => \N__46643\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \N__49522\
        );

    \phase_controller_inst1.start_timer_hc_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__44542\,
            in1 => \N__33366\,
            in2 => \N__33067\,
            in3 => \N__33094\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => 'H',
            sr => \N__49522\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33088\,
            in2 => \_gnd_net_\,
            in3 => \N__33062\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34659\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34918\,
            lcout => \phase_controller_inst1.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46598\,
            in2 => \_gnd_net_\,
            in3 => \N__44618\,
            lcout => \phase_controller_inst1.N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__34957\,
            in1 => \N__34877\,
            in2 => \_gnd_net_\,
            in3 => \N__34850\,
            lcout => \current_shift_inst.timer_s1.N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33295\,
            in2 => \_gnd_net_\,
            in3 => \N__33316\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_13_4_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33268\,
            in3 => \N__33289\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33238\,
            in2 => \_gnd_net_\,
            in3 => \N__33259\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33211\,
            in2 => \_gnd_net_\,
            in3 => \N__33232\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33205\,
            in2 => \_gnd_net_\,
            in3 => \N__33193\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33190\,
            in2 => \_gnd_net_\,
            in3 => \N__33178\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33484\,
            in2 => \_gnd_net_\,
            in3 => \N__33472\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33469\,
            in2 => \_gnd_net_\,
            in3 => \N__33451\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33448\,
            in2 => \_gnd_net_\,
            in3 => \N__33436\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_8\,
            ltout => OPEN,
            carryin => \bfn_13_5_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34993\,
            in2 => \_gnd_net_\,
            in3 => \N__33424\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33421\,
            in2 => \_gnd_net_\,
            in3 => \N__33403\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33400\,
            in2 => \_gnd_net_\,
            in3 => \N__33382\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34753\,
            in2 => \_gnd_net_\,
            in3 => \N__33379\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33727\,
            in2 => \_gnd_net_\,
            in3 => \N__33370\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35036\,
            in2 => \_gnd_net_\,
            in3 => \N__33571\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34746\,
            in2 => \_gnd_net_\,
            in3 => \N__33568\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34140\,
            in2 => \_gnd_net_\,
            in3 => \N__33559\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35486\,
            in2 => \_gnd_net_\,
            in3 => \N__33550\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33545\,
            in2 => \_gnd_net_\,
            in3 => \N__33517\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34979\,
            in2 => \_gnd_net_\,
            in3 => \N__33505\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38057\,
            in2 => \_gnd_net_\,
            in3 => \N__33502\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35340\,
            in2 => \_gnd_net_\,
            in3 => \N__33490\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35078\,
            in2 => \_gnd_net_\,
            in3 => \N__33487\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35207\,
            in2 => \_gnd_net_\,
            in3 => \N__33655\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35307\,
            in3 => \N__33646\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33642\,
            in2 => \_gnd_net_\,
            in3 => \N__33625\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35510\,
            in2 => \_gnd_net_\,
            in3 => \N__33616\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34111\,
            in2 => \_gnd_net_\,
            in3 => \N__33607\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35469\,
            in2 => \_gnd_net_\,
            in3 => \N__33604\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34173\,
            in2 => \_gnd_net_\,
            in3 => \N__33595\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35579\,
            in2 => \_gnd_net_\,
            in3 => \N__33586\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un7_integrator1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__34086\,
            in1 => \N__37946\,
            in2 => \_gnd_net_\,
            in3 => \N__34042\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__37287\,
            in1 => \N__37495\,
            in2 => \N__34027\,
            in3 => \N__37612\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49420\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__37288\,
            in1 => \N__37496\,
            in2 => \N__33979\,
            in3 => \N__37613\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49420\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111110101"
        )
    port map (
            in0 => \N__37493\,
            in1 => \N__37290\,
            in2 => \N__37668\,
            in3 => \N__33967\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49420\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111001110"
        )
    port map (
            in0 => \N__37286\,
            in1 => \N__37494\,
            in2 => \N__33895\,
            in3 => \N__37614\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49420\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111110"
        )
    port map (
            in0 => \N__37492\,
            in1 => \N__37289\,
            in2 => \N__37667\,
            in3 => \N__33883\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49420\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33792\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33743\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33717\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__34139\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37791\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35442\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37792\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34110\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__41634\,
            in1 => \N__38427\,
            in2 => \N__38500\,
            in3 => \N__41808\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49926\,
            ce => \N__36763\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__41807\,
            in1 => \N__38522\,
            in2 => \N__38431\,
            in3 => \N__41637\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49926\,
            ce => \N__36763\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__41633\,
            in1 => \N__38426\,
            in2 => \N__38572\,
            in3 => \N__41805\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49926\,
            ce => \N__36763\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__41635\,
            in1 => \N__41809\,
            in2 => \N__41449\,
            in3 => \N__38428\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49926\,
            ce => \N__36763\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__41806\,
            in1 => \N__38547\,
            in2 => \N__38430\,
            in3 => \N__41636\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49926\,
            ce => \N__36763\,
            sr => \N__49432\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36817\,
            in2 => \_gnd_net_\,
            in3 => \N__36838\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37050\,
            in2 => \_gnd_net_\,
            in3 => \N__36796\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__49583\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34172\,
            in2 => \_gnd_net_\,
            in3 => \N__37833\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__38769\,
            in1 => \N__41781\,
            in2 => \N__40642\,
            in3 => \N__38851\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49915\,
            ce => \N__36761\,
            sr => \N__49449\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__35733\,
            in1 => \N__38844\,
            in2 => \N__38791\,
            in3 => \N__40692\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49915\,
            ce => \N__36761\,
            sr => \N__49449\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__38768\,
            in1 => \N__41779\,
            in2 => \N__41104\,
            in3 => \N__38850\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49915\,
            ce => \N__36761\,
            sr => \N__49449\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__35715\,
            in1 => \N__38776\,
            in2 => \_gnd_net_\,
            in3 => \N__41777\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49915\,
            ce => \N__36761\,
            sr => \N__49449\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__41780\,
            in1 => \N__38845\,
            in2 => \N__41143\,
            in3 => \N__38770\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49915\,
            ce => \N__36761\,
            sr => \N__49449\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__41778\,
            in1 => \N__35676\,
            in2 => \_gnd_net_\,
            in3 => \N__38771\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49915\,
            ce => \N__36761\,
            sr => \N__49449\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35752\,
            in2 => \N__34153\,
            in3 => \N__36074\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36049\,
            in1 => \N__35746\,
            in2 => \N__34309\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34300\,
            in2 => \N__34294\,
            in3 => \N__36022\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34282\,
            in2 => \N__34276\,
            in3 => \N__36004\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34267\,
            in2 => \N__34261\,
            in3 => \N__35986\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34249\,
            in2 => \N__34243\,
            in3 => \N__36391\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36370\,
            in1 => \N__34225\,
            in2 => \N__34234\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34210\,
            in2 => \N__34219\,
            in3 => \N__36352\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36334\,
            in1 => \N__34204\,
            in2 => \N__35557\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34402\,
            in2 => \N__34414\,
            in3 => \N__36316\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34396\,
            in2 => \N__34387\,
            in3 => \N__36298\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34375\,
            in2 => \N__34366\,
            in3 => \N__36274\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34357\,
            in2 => \N__34348\,
            in3 => \N__36256\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36556\,
            in1 => \N__34336\,
            in2 => \N__34327\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35542\,
            in2 => \N__34318\,
            in3 => \N__36538\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35890\,
            in2 => \N__35530\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35941\,
            in2 => \N__35968\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36985\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36943\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36904\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36865\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34438\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34429\,
            in2 => \N__37057\,
            in3 => \N__34420\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34417\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__42267\,
            in1 => \N__34608\,
            in2 => \N__42220\,
            in3 => \N__34482\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49894\,
            ce => \N__49122\,
            sr => \N__49479\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39340\,
            in1 => \N__39357\,
            in2 => \N__45631\,
            in3 => \N__39372\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__39358\,
            in1 => \N__45560\,
            in2 => \N__45936\,
            in3 => \N__34506\,
            lcout => \elapsed_time_ns_1_RNIPKKEE1_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__45929\,
            in1 => \N__39373\,
            in2 => \N__45562\,
            in3 => \N__38312\,
            lcout => \elapsed_time_ns_1_RNIOJKEE1_0_7\,
            ltout => \elapsed_time_ns_1_RNIOJKEE1_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__45959\,
            in1 => \N__34505\,
            in2 => \N__34492\,
            in3 => \N__45786\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46746\,
            in2 => \N__34489\,
            in3 => \N__45705\,
            lcout => \phase_controller_inst1.stoper_hc.N_330\,
            ltout => \phase_controller_inst1.stoper_hc.N_330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__45960\,
            in1 => \N__47084\,
            in2 => \N__34486\,
            in3 => \N__42212\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49888\,
            ce => \N__49109\,
            sr => \N__49486\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__46747\,
            in1 => \N__47083\,
            in2 => \N__34459\,
            in3 => \N__34471\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100110011"
        )
    port map (
            in0 => \N__34455\,
            in1 => \N__34572\,
            in2 => \N__34607\,
            in3 => \N__34470\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__34552\,
            in1 => \N__45937\,
            in2 => \N__34576\,
            in3 => \N__45548\,
            lcout => \elapsed_time_ns_1_RNIJEKEE1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__45588\,
            in1 => \N__46874\,
            in2 => \N__45730\,
            in3 => \N__37021\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2\,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34561\,
            in1 => \N__34454\,
            in2 => \N__34441\,
            in3 => \N__46800\,
            lcout => \phase_controller_inst1.stoper_hc.N_310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34597\,
            in2 => \_gnd_net_\,
            in3 => \N__34571\,
            lcout => \phase_controller_inst1.stoper_hc.N_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46048\,
            in2 => \_gnd_net_\,
            in3 => \N__42331\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__39223\,
            in1 => \N__39240\,
            in2 => \N__34555\,
            in3 => \N__34551\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39759\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49881\,
            ce => \N__39447\,
            sr => \N__49492\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__46886\,
            in1 => \N__45589\,
            in2 => \_gnd_net_\,
            in3 => \N__45787\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010000"
        )
    port map (
            in0 => \N__45731\,
            in1 => \N__46812\,
            in2 => \N__34543\,
            in3 => \N__45668\,
            lcout => \phase_controller_inst1.stoper_hc.N_328\,
            ltout => \phase_controller_inst1.stoper_hc.N_328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47078\,
            in2 => \N__34540\,
            in3 => \N__34533\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011111110"
        )
    port map (
            in0 => \N__34532\,
            in1 => \N__45561\,
            in2 => \N__45379\,
            in3 => \N__39463\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34537\,
            in3 => \N__46024\,
            lcout => \elapsed_time_ns_1_RNIP93CP1_0_1\,
            ltout => \elapsed_time_ns_1_RNIP93CP1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__42271\,
            in1 => \N__34734\,
            in2 => \N__34723\,
            in3 => \N__34719\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49874\,
            ce => \N__49110\,
            sr => \N__49501\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__34701\,
            in1 => \N__42193\,
            in2 => \N__42285\,
            in3 => \N__47079\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49874\,
            ce => \N__49110\,
            sr => \N__49501\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__42192\,
            in1 => \N__42272\,
            in2 => \N__47105\,
            in3 => \N__39307\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49874\,
            ce => \N__49110\,
            sr => \N__49501\
        );

    \phase_controller_inst2.state_3_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__41246\,
            in1 => \N__34672\,
            in2 => \N__41227\,
            in3 => \N__35818\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49869\,
            ce => 'H',
            sr => \N__49507\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__47111\,
            in1 => \N__46801\,
            in2 => \N__45736\,
            in3 => \N__45672\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49864\,
            ce => \N__43143\,
            sr => \N__49513\
        );

    \phase_controller_inst1.state_3_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__38257\,
            in1 => \N__34671\,
            in2 => \N__38296\,
            in3 => \N__44490\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49859\,
            ce => 'H',
            sr => \N__49517\
        );

    \phase_controller_inst1.state_0_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__44602\,
            in1 => \N__34660\,
            in2 => \N__46656\,
            in3 => \N__34920\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49857\,
            ce => 'H',
            sr => \N__49523\
        );

    \phase_controller_inst1.T45_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__38254\,
            in1 => \N__34620\,
            in2 => \_gnd_net_\,
            in3 => \N__34919\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49857\,
            ce => 'H',
            sr => \N__49523\
        );

    \current_shift_inst.stop_timer_s1_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__38259\,
            in1 => \N__34935\,
            in2 => \N__34963\,
            in3 => \N__34851\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49853\,
            ce => 'H',
            sr => \N__49525\
        );

    \current_shift_inst.timer_s1.running_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__34852\,
            in1 => \N__34962\,
            in2 => \_gnd_net_\,
            in3 => \N__34878\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49853\,
            ce => 'H',
            sr => \N__49525\
        );

    \current_shift_inst.start_timer_s1_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__34934\,
            in1 => \N__34961\,
            in2 => \_gnd_net_\,
            in3 => \N__38258\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49853\,
            ce => 'H',
            sr => \N__49525\
        );

    \phase_controller_inst1.S1_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38260\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49853\,
            ce => 'H',
            sr => \N__49525\
        );

    \phase_controller_inst1.T23_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__34890\,
            in1 => \N__46664\,
            in2 => \_gnd_net_\,
            in3 => \N__34921\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49853\,
            ce => 'H',
            sr => \N__49525\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34873\,
            in2 => \_gnd_net_\,
            in3 => \N__34849\,
            lcout => \current_shift_inst.timer_s1.N_166_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46663\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49850\,
            ce => 'H',
            sr => \N__49532\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__37666\,
            in1 => \N__37323\,
            in2 => \_gnd_net_\,
            in3 => \N__34813\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49964\,
            ce => 'H',
            sr => \N__49405\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35190\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__34747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37976\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110101"
        )
    port map (
            in0 => \N__37979\,
            in1 => \N__35283\,
            in2 => \N__35239\,
            in3 => \N__35236\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__35080\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37977\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__35211\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37978\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__37082\,
            in1 => \N__37950\,
            in2 => \N__35191\,
            in3 => \N__35152\,
            lcout => \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111001111"
        )
    port map (
            in0 => \N__35131\,
            in1 => \N__35079\,
            in2 => \N__37975\,
            in3 => \N__35062\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__35040\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37947\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35019\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__38059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37949\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__34983\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37948\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__35514\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37934\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__35490\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37933\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35470\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28\,
            ltout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111110011"
        )
    port map (
            in0 => \N__35458\,
            in1 => \N__37936\,
            in2 => \N__35407\,
            in3 => \N__35404\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35382\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__35339\,
            in1 => \N__37937\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38004\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37938\,
            in2 => \_gnd_net_\,
            in3 => \N__35306\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35651\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38086\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37939\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35583\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__41319\,
            in1 => \N__38467\,
            in2 => \_gnd_net_\,
            in3 => \N__35776\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011100"
        )
    port map (
            in0 => \N__41594\,
            in1 => \N__41761\,
            in2 => \N__35563\,
            in3 => \N__38659\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__41320\,
            in1 => \N__41596\,
            in2 => \N__35560\,
            in3 => \N__38429\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49939\,
            ce => \N__36754\,
            sr => \N__49421\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__38468\,
            in1 => \N__41763\,
            in2 => \N__41630\,
            in3 => \N__38692\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49939\,
            ce => \N__36754\,
            sr => \N__49421\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__41762\,
            in1 => \N__41595\,
            in2 => \_gnd_net_\,
            in3 => \N__41968\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49939\,
            ce => \N__36754\,
            sr => \N__49421\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__35908\,
            in1 => \N__35922\,
            in2 => \N__36517\,
            in3 => \N__36477\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__41023\,
            in1 => \N__44053\,
            in2 => \N__40816\,
            in3 => \N__38524\,
            lcout => \elapsed_time_ns_1_RNIR9HF91_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__38548\,
            in1 => \N__44101\,
            in2 => \N__40818\,
            in3 => \N__41024\,
            lcout => \elapsed_time_ns_1_RNIQ8HF91_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__41025\,
            in1 => \N__35714\,
            in2 => \N__40817\,
            in3 => \N__47275\,
            lcout => \elapsed_time_ns_1_RNIFJ2591_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__41444\,
            in1 => \N__38684\,
            in2 => \_gnd_net_\,
            in3 => \N__38469\,
            lcout => \phase_controller_inst1.stoper_tr.N_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__41022\,
            in1 => \N__44011\,
            in2 => \N__40815\,
            in3 => \N__38499\,
            lcout => \elapsed_time_ns_1_RNISAHF91_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__35675\,
            in1 => \N__41054\,
            in2 => \N__47302\,
            in3 => \N__40822\,
            lcout => \elapsed_time_ns_1_RNIGK2591_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__41770\,
            in1 => \N__38622\,
            in2 => \N__38643\,
            in3 => \N__41625\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__40821\,
            in1 => \N__38564\,
            in2 => \N__41061\,
            in3 => \N__43480\,
            lcout => \elapsed_time_ns_1_RNIP7HF91_0_10\,
            ltout => \elapsed_time_ns_1_RNIP7HF91_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38494\,
            in1 => \N__38521\,
            in2 => \N__35722\,
            in3 => \N__38545\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__35707\,
            in1 => \N__40634\,
            in2 => \N__35686\,
            in3 => \N__35674\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__38470\,
            in1 => \_gnd_net_\,
            in2 => \N__35779\,
            in3 => \N__41624\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__38623\,
            in1 => \N__40685\,
            in2 => \N__38644\,
            in3 => \N__38608\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__38472\,
            in1 => \N__41310\,
            in2 => \_gnd_net_\,
            in3 => \N__41432\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__41433\,
            in1 => \N__41311\,
            in2 => \_gnd_net_\,
            in3 => \N__35772\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__38683\,
            in1 => \N__38473\,
            in2 => \N__35761\,
            in3 => \N__41626\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111010"
        )
    port map (
            in0 => \N__41698\,
            in1 => \_gnd_net_\,
            in2 => \N__35758\,
            in3 => \N__38910\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__38911\,
            in1 => \N__38896\,
            in2 => \N__35755\,
            in3 => \N__38849\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49921\,
            ce => \N__36750\,
            sr => \N__49439\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__41699\,
            in1 => \N__38874\,
            in2 => \N__38856\,
            in3 => \N__38780\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49921\,
            ce => \N__36750\,
            sr => \N__49439\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__45354\,
            in1 => \N__41875\,
            in2 => \N__41062\,
            in3 => \N__47173\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__41751\,
            in1 => \N__41874\,
            in2 => \_gnd_net_\,
            in3 => \N__41629\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49916\,
            ce => \N__36762\,
            sr => \N__49450\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__36420\,
            in1 => \N__35931\,
            in2 => \N__36448\,
            in3 => \N__35949\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__35932\,
            in1 => \N__36447\,
            in2 => \N__35953\,
            in3 => \N__36421\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__41627\,
            in1 => \N__41750\,
            in2 => \_gnd_net_\,
            in3 => \N__41503\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49916\,
            ce => \N__36762\,
            sr => \N__49450\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__41749\,
            in1 => \N__41923\,
            in2 => \_gnd_net_\,
            in3 => \N__41628\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49916\,
            ce => \N__36762\,
            sr => \N__49450\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__36478\,
            in1 => \N__35923\,
            in2 => \N__36516\,
            in3 => \N__35904\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__35883\,
            in1 => \N__41197\,
            in2 => \N__46201\,
            in3 => \N__35843\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__35817\,
            in1 => \N__36170\,
            in2 => \N__35797\,
            in3 => \N__44553\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49457\
        );

    \phase_controller_inst2.stoper_tr.running_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011111010"
        )
    port map (
            in0 => \N__36190\,
            in1 => \N__35793\,
            in2 => \N__36142\,
            in3 => \N__36224\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49457\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111011101"
        )
    port map (
            in0 => \N__36223\,
            in1 => \N__37043\,
            in2 => \N__36795\,
            in3 => \N__36238\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36232\,
            in3 => \N__36125\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__36222\,
            in1 => \N__36189\,
            in2 => \_gnd_net_\,
            in3 => \N__36163\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => \phase_controller_inst2.stoper_tr.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36109\,
            in3 => \N__36099\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36088\,
            in2 => \N__36082\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36743\,
            in1 => \N__36048\,
            in2 => \_gnd_net_\,
            in3 => \N__36034\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49464\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__36747\,
            in1 => \N__36021\,
            in2 => \N__36031\,
            in3 => \N__36007\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49464\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36744\,
            in1 => \N__36003\,
            in2 => \_gnd_net_\,
            in3 => \N__35989\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49464\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36748\,
            in1 => \N__35985\,
            in2 => \_gnd_net_\,
            in3 => \N__35971\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49464\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36745\,
            in1 => \N__36387\,
            in2 => \_gnd_net_\,
            in3 => \N__36373\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49464\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36749\,
            in1 => \N__36369\,
            in2 => \_gnd_net_\,
            in3 => \N__36355\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49464\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36746\,
            in1 => \N__36351\,
            in2 => \_gnd_net_\,
            in3 => \N__36337\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49906\,
            ce => 'H',
            sr => \N__49464\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36729\,
            in1 => \N__36333\,
            in2 => \_gnd_net_\,
            in3 => \N__36319\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36696\,
            in1 => \N__36315\,
            in2 => \_gnd_net_\,
            in3 => \N__36301\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36726\,
            in1 => \N__36291\,
            in2 => \_gnd_net_\,
            in3 => \N__36277\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36697\,
            in1 => \N__36273\,
            in2 => \_gnd_net_\,
            in3 => \N__36259\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36727\,
            in1 => \N__36255\,
            in2 => \_gnd_net_\,
            in3 => \N__36241\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36698\,
            in1 => \N__36555\,
            in2 => \_gnd_net_\,
            in3 => \N__36541\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36728\,
            in1 => \N__36534\,
            in2 => \_gnd_net_\,
            in3 => \N__36520\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36699\,
            in1 => \N__36500\,
            in2 => \_gnd_net_\,
            in3 => \N__36481\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49900\,
            ce => 'H',
            sr => \N__49471\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36692\,
            in1 => \N__36473\,
            in2 => \_gnd_net_\,
            in3 => \N__36451\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49895\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36722\,
            in1 => \N__36438\,
            in2 => \_gnd_net_\,
            in3 => \N__36424\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49895\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36693\,
            in1 => \N__36419\,
            in2 => \_gnd_net_\,
            in3 => \N__36403\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49895\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36723\,
            in1 => \N__36999\,
            in2 => \_gnd_net_\,
            in3 => \N__36400\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49895\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36694\,
            in1 => \N__37014\,
            in2 => \_gnd_net_\,
            in3 => \N__36397\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49895\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36724\,
            in1 => \N__36957\,
            in2 => \_gnd_net_\,
            in3 => \N__36394\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49895\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36695\,
            in1 => \N__36972\,
            in2 => \_gnd_net_\,
            in3 => \N__36853\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49895\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36725\,
            in1 => \N__36930\,
            in2 => \_gnd_net_\,
            in3 => \N__36850\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49895\,
            ce => 'H',
            sr => \N__49480\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36688\,
            in1 => \N__36916\,
            in2 => \_gnd_net_\,
            in3 => \N__36847\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49487\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36719\,
            in1 => \N__36879\,
            in2 => \_gnd_net_\,
            in3 => \N__36844\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49487\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36689\,
            in1 => \N__36892\,
            in2 => \_gnd_net_\,
            in3 => \N__36841\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49487\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36720\,
            in1 => \N__36834\,
            in2 => \_gnd_net_\,
            in3 => \N__36820\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49487\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36690\,
            in1 => \N__36813\,
            in2 => \_gnd_net_\,
            in3 => \N__36799\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49487\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36721\,
            in1 => \N__36788\,
            in2 => \_gnd_net_\,
            in3 => \N__36766\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49487\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36691\,
            in1 => \N__37042\,
            in2 => \_gnd_net_\,
            in3 => \N__37060\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49487\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48286\,
            in2 => \_gnd_net_\,
            in3 => \N__47968\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47992\,
            in2 => \_gnd_net_\,
            in3 => \N__48013\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__45208\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46023\,
            lcout => \elapsed_time_ns_1_RNI1I3CP1_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__42775\,
            in1 => \N__42646\,
            in2 => \_gnd_net_\,
            in3 => \N__39268\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__37015\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37000\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36973\,
            in2 => \_gnd_net_\,
            in3 => \N__36958\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__36931\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36915\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__36891\,
            in1 => \_gnd_net_\,
            in2 => \N__36880\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__47106\,
            in1 => \N__38322\,
            in2 => \_gnd_net_\,
            in3 => \N__42205\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49875\,
            ce => \N__49121\,
            sr => \N__49502\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__47107\,
            in1 => \N__45757\,
            in2 => \N__45602\,
            in3 => \N__46826\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49875\,
            ce => \N__49121\,
            sr => \N__49502\
        );

    \phase_controller_inst1.state_2_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__38294\,
            in1 => \N__46587\,
            in2 => \N__44640\,
            in3 => \N__38255\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49865\,
            ce => 'H',
            sr => \N__49514\
        );

    \phase_controller_inst1.T01_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__38202\,
            in1 => \N__38256\,
            in2 => \_gnd_net_\,
            in3 => \N__46588\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49860\,
            ce => 'H',
            sr => \N__49518\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011111110"
        )
    port map (
            in0 => \N__37713\,
            in1 => \N__37498\,
            in2 => \N__37326\,
            in3 => \N__38191\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49965\,
            ce => 'H',
            sr => \N__49406\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000111110101"
        )
    port map (
            in0 => \N__37501\,
            in1 => \N__37284\,
            in2 => \N__37714\,
            in3 => \N__38122\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49960\,
            ce => 'H',
            sr => \N__49408\
        );

    \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110101111"
        )
    port map (
            in0 => \N__38058\,
            in1 => \N__38035\,
            in2 => \N__37984\,
            in3 => \N__37738\,
            lcout => \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000110111011"
        )
    port map (
            in0 => \N__37709\,
            in1 => \N__37497\,
            in2 => \N__37327\,
            in3 => \N__37123\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49954\,
            ce => 'H',
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__40972\,
            in1 => \N__38374\,
            in2 => \N__44206\,
            in3 => \N__40779\,
            lcout => \elapsed_time_ns_1_RNIVEIF91_0_25\,
            ltout => \elapsed_time_ns_1_RNIVEIF91_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38364\,
            in1 => \N__38352\,
            in2 => \N__38368\,
            in3 => \N__38583\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__40973\,
            in1 => \N__38365\,
            in2 => \N__44857\,
            in3 => \N__40780\,
            lcout => \elapsed_time_ns_1_RNI2IIF91_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__40974\,
            in1 => \N__44914\,
            in2 => \N__38356\,
            in3 => \N__40781\,
            lcout => \elapsed_time_ns_1_RNI1HIF91_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40255\,
            in1 => \N__38344\,
            in2 => \N__40597\,
            in3 => \N__38331\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_19_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__49580\,
            in1 => \N__41173\,
            in2 => \N__47455\,
            in3 => \N__45290\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111100"
        )
    port map (
            in0 => \N__44695\,
            in1 => \N__49581\,
            in2 => \N__38338\,
            in3 => \N__47719\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31\,
            ltout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__44377\,
            in1 => \N__41007\,
            in2 => \N__38335\,
            in3 => \N__40279\,
            lcout => \elapsed_time_ns_1_RNIRAIF91_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__38332\,
            in1 => \N__44338\,
            in2 => \N__41049\,
            in3 => \N__40785\,
            lcout => \elapsed_time_ns_1_RNISBIF91_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__41395\,
            in1 => \N__44694\,
            in2 => \_gnd_net_\,
            in3 => \N__41380\,
            lcout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i\,
            ltout => \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__38584\,
            in1 => \N__44161\,
            in2 => \N__38587\,
            in3 => \N__40784\,
            lcout => \elapsed_time_ns_1_RNI0GIF91_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__41775\,
            in1 => \N__41448\,
            in2 => \N__41623\,
            in3 => \N__38419\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => \N__50322\,
            sr => \N__49422\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__38414\,
            in1 => \N__41568\,
            in2 => \N__38571\,
            in3 => \N__41771\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => \N__50322\,
            sr => \N__49422\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__41772\,
            in1 => \N__38417\,
            in2 => \N__41621\,
            in3 => \N__38546\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => \N__50322\,
            sr => \N__49422\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__38415\,
            in1 => \N__38523\,
            in2 => \N__41632\,
            in3 => \N__41773\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => \N__50322\,
            sr => \N__49422\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__41774\,
            in1 => \N__38418\,
            in2 => \N__41622\,
            in3 => \N__38495\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => \N__50322\,
            sr => \N__49422\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__43930\,
            in1 => \N__38471\,
            in2 => \N__41050\,
            in3 => \N__40788\,
            lcout => \elapsed_time_ns_1_RNIUCHF91_0_15\,
            ltout => \elapsed_time_ns_1_RNIUCHF91_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__41776\,
            in1 => \N__41600\,
            in2 => \N__38434\,
            in3 => \N__38688\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => \N__50322\,
            sr => \N__49422\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__38416\,
            in1 => \N__41317\,
            in2 => \N__41631\,
            in3 => \N__38380\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => \N__50322\,
            sr => \N__49422\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__41955\,
            in1 => \N__41911\,
            in2 => \N__41498\,
            in3 => \N__41861\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__38607\,
            in1 => \N__41055\,
            in2 => \N__47368\,
            in3 => \N__40819\,
            lcout => \elapsed_time_ns_1_RNIAE2591_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_7_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__40856\,
            in1 => \N__41168\,
            in2 => \_gnd_net_\,
            in3 => \N__40835\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__47311\,
            in1 => \_gnd_net_\,
            in2 => \N__38662\,
            in3 => \N__47711\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__41956\,
            in1 => \N__41068\,
            in2 => \N__41918\,
            in3 => \N__38655\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__38593\,
            in1 => \N__41593\,
            in2 => \N__38626\,
            in3 => \N__38621\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__40674\,
            in1 => \N__38606\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_19_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__41169\,
            in1 => \N__40857\,
            in2 => \N__40840\,
            in3 => \N__47451\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101110"
        )
    port map (
            in0 => \N__45348\,
            in1 => \N__41056\,
            in2 => \N__47332\,
            in3 => \N__38909\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38914\,
            in3 => \N__41365\,
            lcout => \elapsed_time_ns_1_RNII6NQL1_0_1\,
            ltout => \elapsed_time_ns_1_RNII6NQL1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__38895\,
            in1 => \N__38839\,
            in2 => \N__38884\,
            in3 => \N__38881\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49927\,
            ce => \N__50323\,
            sr => \N__49433\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__38838\,
            in1 => \N__41769\,
            in2 => \N__38790\,
            in3 => \N__40630\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49927\,
            ce => \N__50323\,
            sr => \N__49433\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__41764\,
            in1 => \N__44693\,
            in2 => \N__41060\,
            in3 => \N__40820\,
            lcout => \elapsed_time_ns_1_RNISCJF91_0_31\,
            ltout => \elapsed_time_ns_1_RNISCJF91_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__38837\,
            in1 => \N__38875\,
            in2 => \N__38863\,
            in3 => \N__38781\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49927\,
            ce => \N__50323\,
            sr => \N__49433\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__41100\,
            in1 => \N__38772\,
            in2 => \N__41802\,
            in3 => \N__38843\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49927\,
            ce => \N__50323\,
            sr => \N__49433\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__41138\,
            in1 => \N__41768\,
            in2 => \N__38855\,
            in3 => \N__38782\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49927\,
            ce => \N__50323\,
            sr => \N__49433\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38713\,
            in2 => \N__38722\,
            in3 => \N__47669\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38698\,
            in2 => \N__38707\,
            in3 => \N__47656\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__47623\,
            in1 => \N__39061\,
            in2 => \N__39049\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__47605\,
            in1 => \N__39040\,
            in2 => \N__39034\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39025\,
            in2 => \N__39019\,
            in3 => \N__47584\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39010\,
            in2 => \N__39004\,
            in3 => \N__47566\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38992\,
            in2 => \N__38980\,
            in3 => \N__47548\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__47527\,
            in1 => \N__38971\,
            in2 => \N__38959\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38950\,
            in2 => \N__38941\,
            in3 => \N__47941\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38932\,
            in2 => \N__38923\,
            in3 => \N__47923\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__47905\,
            in1 => \N__39142\,
            in2 => \N__39154\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39136\,
            in2 => \N__39127\,
            in3 => \N__47887\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39118\,
            in2 => \N__39109\,
            in3 => \N__47869\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39100\,
            in2 => \N__39091\,
            in3 => \N__47851\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39079\,
            in2 => \N__39070\,
            in3 => \N__47833\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41974\,
            in2 => \N__41989\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41815\,
            in2 => \N__41839\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48847\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39196\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39184\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45025\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45037\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44953\,
            in2 => \N__48178\,
            in3 => \N__39172\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39169\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42045\,
            in1 => \N__39249\,
            in2 => \N__39166\,
            in3 => \N__39258\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__45861\,
            in1 => \N__39489\,
            in2 => \N__45511\,
            in3 => \N__39165\,
            lcout => \elapsed_time_ns_1_RNI4HV8E1_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__45459\,
            in1 => \N__45868\,
            in2 => \N__42475\,
            in3 => \N__45169\,
            lcout => \elapsed_time_ns_1_RNI8KU8E1_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__45860\,
            in1 => \N__45455\,
            in2 => \N__39296\,
            in3 => \N__39219\,
            lcout => \elapsed_time_ns_1_RNILGKEE1_0_4\,
            ltout => \elapsed_time_ns_1_RNILGKEE1_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42302\,
            in1 => \N__42954\,
            in2 => \N__39271\,
            in3 => \N__43375\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__39259\,
            in1 => \N__42034\,
            in2 => \N__45905\,
            in3 => \N__45458\,
            lcout => \elapsed_time_ns_1_RNI4GU8E1_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__45456\,
            in1 => \N__43297\,
            in2 => \N__45927\,
            in3 => \N__39339\,
            lcout => \elapsed_time_ns_1_RNI2DT8E1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__39250\,
            in1 => \N__39517\,
            in2 => \N__45904\,
            in3 => \N__45457\,
            lcout => \elapsed_time_ns_1_RNICOU8E1_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39723\,
            in2 => \N__39430\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49901\,
            ce => \N__39451\,
            sr => \N__49472\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39702\,
            in2 => \N__39760\,
            in3 => \N__39205\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49901\,
            ce => \N__39451\,
            sr => \N__49472\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39724\,
            in2 => \N__39679\,
            in3 => \N__39202\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49901\,
            ce => \N__39451\,
            sr => \N__49472\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39703\,
            in2 => \N__39651\,
            in3 => \N__39199\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49901\,
            ce => \N__39451\,
            sr => \N__49472\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39678\,
            in2 => \N__39621\,
            in3 => \N__39361\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49901\,
            ce => \N__39451\,
            sr => \N__49472\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39588\,
            in2 => \N__39652\,
            in3 => \N__39346\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49901\,
            ce => \N__39451\,
            sr => \N__49472\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39555\,
            in2 => \N__39622\,
            in3 => \N__39343\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49901\,
            ce => \N__39451\,
            sr => \N__49472\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39987\,
            in2 => \N__39592\,
            in3 => \N__39325\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49901\,
            ce => \N__39451\,
            sr => \N__49472\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39960\,
            in2 => \N__39562\,
            in3 => \N__39322\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49896\,
            ce => \N__39450\,
            sr => \N__49481\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39936\,
            in2 => \N__39991\,
            in3 => \N__39319\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49896\,
            ce => \N__39450\,
            sr => \N__49481\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39961\,
            in2 => \N__39912\,
            in3 => \N__39316\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49896\,
            ce => \N__39450\,
            sr => \N__49481\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39937\,
            in2 => \N__39882\,
            in3 => \N__39313\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49896\,
            ce => \N__39450\,
            sr => \N__49481\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39849\,
            in2 => \N__39913\,
            in3 => \N__39310\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49896\,
            ce => \N__39450\,
            sr => \N__49481\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39819\,
            in2 => \N__39883\,
            in3 => \N__39400\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49896\,
            ce => \N__39450\,
            sr => \N__49481\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39789\,
            in2 => \N__39853\,
            in3 => \N__39397\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49896\,
            ce => \N__39450\,
            sr => \N__49481\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40239\,
            in2 => \N__39823\,
            in3 => \N__39394\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49896\,
            ce => \N__39450\,
            sr => \N__49481\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40209\,
            in2 => \N__39793\,
            in3 => \N__39391\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49890\,
            ce => \N__39449\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40243\,
            in2 => \N__40182\,
            in3 => \N__39388\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49890\,
            ce => \N__39449\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40155\,
            in2 => \N__40213\,
            in3 => \N__39385\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49890\,
            ce => \N__39449\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40131\,
            in2 => \N__40183\,
            in3 => \N__39382\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49890\,
            ce => \N__39449\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40156\,
            in2 => \N__40107\,
            in3 => \N__39379\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49890\,
            ce => \N__39449\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40077\,
            in2 => \N__40135\,
            in3 => \N__39376\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49890\,
            ce => \N__39449\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40050\,
            in2 => \N__40108\,
            in3 => \N__39529\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49890\,
            ce => \N__39449\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40078\,
            in2 => \N__40023\,
            in3 => \N__39526\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49890\,
            ce => \N__39449\,
            sr => \N__49488\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40551\,
            in2 => \N__40057\,
            in3 => \N__39523\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49882\,
            ce => \N__39448\,
            sr => \N__49493\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40024\,
            in2 => \N__40530\,
            in3 => \N__39520\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49882\,
            ce => \N__39448\,
            sr => \N__49493\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40552\,
            in2 => \N__40504\,
            in3 => \N__39496\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49882\,
            ce => \N__39448\,
            sr => \N__49493\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40342\,
            in2 => \N__40531\,
            in3 => \N__39469\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49882\,
            ce => \N__39448\,
            sr => \N__49493\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39466\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49882\,
            ce => \N__39448\,
            sr => \N__49493\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39423\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49882\,
            ce => \N__39448\,
            sr => \N__49493\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40476\,
            in1 => \N__39422\,
            in2 => \_gnd_net_\,
            in3 => \N__39403\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__49876\,
            ce => \N__40318\,
            sr => \N__49503\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40480\,
            in1 => \N__39746\,
            in2 => \_gnd_net_\,
            in3 => \N__39727\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__49876\,
            ce => \N__40318\,
            sr => \N__49503\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40477\,
            in1 => \N__39722\,
            in2 => \_gnd_net_\,
            in3 => \N__39706\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__49876\,
            ce => \N__40318\,
            sr => \N__49503\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40481\,
            in1 => \N__39696\,
            in2 => \_gnd_net_\,
            in3 => \N__39682\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__49876\,
            ce => \N__40318\,
            sr => \N__49503\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40478\,
            in1 => \N__39674\,
            in2 => \_gnd_net_\,
            in3 => \N__39655\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__49876\,
            ce => \N__40318\,
            sr => \N__49503\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40482\,
            in1 => \N__39639\,
            in2 => \_gnd_net_\,
            in3 => \N__39625\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__49876\,
            ce => \N__40318\,
            sr => \N__49503\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40479\,
            in1 => \N__39609\,
            in2 => \_gnd_net_\,
            in3 => \N__39595\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__49876\,
            ce => \N__40318\,
            sr => \N__49503\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40483\,
            in1 => \N__39581\,
            in2 => \_gnd_net_\,
            in3 => \N__39565\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__49876\,
            ce => \N__40318\,
            sr => \N__49503\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40404\,
            in1 => \N__39554\,
            in2 => \_gnd_net_\,
            in3 => \N__39532\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__49870\,
            ce => \N__40326\,
            sr => \N__49508\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40443\,
            in1 => \N__39980\,
            in2 => \_gnd_net_\,
            in3 => \N__39964\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__49870\,
            ce => \N__40326\,
            sr => \N__49508\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40401\,
            in1 => \N__39954\,
            in2 => \_gnd_net_\,
            in3 => \N__39940\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__49870\,
            ce => \N__40326\,
            sr => \N__49508\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40440\,
            in1 => \N__39930\,
            in2 => \_gnd_net_\,
            in3 => \N__39916\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__49870\,
            ce => \N__40326\,
            sr => \N__49508\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40402\,
            in1 => \N__39900\,
            in2 => \_gnd_net_\,
            in3 => \N__39886\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__49870\,
            ce => \N__40326\,
            sr => \N__49508\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40441\,
            in1 => \N__39870\,
            in2 => \_gnd_net_\,
            in3 => \N__39856\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__49870\,
            ce => \N__40326\,
            sr => \N__49508\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40403\,
            in1 => \N__39842\,
            in2 => \_gnd_net_\,
            in3 => \N__39826\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__49870\,
            ce => \N__40326\,
            sr => \N__49508\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40442\,
            in1 => \N__39812\,
            in2 => \_gnd_net_\,
            in3 => \N__39796\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__49870\,
            ce => \N__40326\,
            sr => \N__49508\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40457\,
            in1 => \N__39782\,
            in2 => \_gnd_net_\,
            in3 => \N__39763\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__49866\,
            ce => \N__40325\,
            sr => \N__49515\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40453\,
            in1 => \N__40238\,
            in2 => \_gnd_net_\,
            in3 => \N__40216\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__49866\,
            ce => \N__40325\,
            sr => \N__49515\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40458\,
            in1 => \N__40202\,
            in2 => \_gnd_net_\,
            in3 => \N__40186\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__49866\,
            ce => \N__40325\,
            sr => \N__49515\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40454\,
            in1 => \N__40175\,
            in2 => \_gnd_net_\,
            in3 => \N__40159\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__49866\,
            ce => \N__40325\,
            sr => \N__49515\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40459\,
            in1 => \N__40154\,
            in2 => \_gnd_net_\,
            in3 => \N__40138\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__49866\,
            ce => \N__40325\,
            sr => \N__49515\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40455\,
            in1 => \N__40130\,
            in2 => \_gnd_net_\,
            in3 => \N__40111\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__49866\,
            ce => \N__40325\,
            sr => \N__49515\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40460\,
            in1 => \N__40095\,
            in2 => \_gnd_net_\,
            in3 => \N__40081\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__49866\,
            ce => \N__40325\,
            sr => \N__49515\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40456\,
            in1 => \N__40076\,
            in2 => \_gnd_net_\,
            in3 => \N__40060\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__49866\,
            ce => \N__40325\,
            sr => \N__49515\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40461\,
            in1 => \N__40049\,
            in2 => \_gnd_net_\,
            in3 => \N__40027\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__49861\,
            ce => \N__40327\,
            sr => \N__49519\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40465\,
            in1 => \N__40016\,
            in2 => \_gnd_net_\,
            in3 => \N__39994\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__49861\,
            ce => \N__40327\,
            sr => \N__49519\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40462\,
            in1 => \N__40550\,
            in2 => \_gnd_net_\,
            in3 => \N__40534\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__49861\,
            ce => \N__40327\,
            sr => \N__49519\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40466\,
            in1 => \N__40523\,
            in2 => \_gnd_net_\,
            in3 => \N__40507\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__49861\,
            ce => \N__40327\,
            sr => \N__49519\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__40463\,
            in1 => \N__40500\,
            in2 => \_gnd_net_\,
            in3 => \N__40486\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__49861\,
            ce => \N__40327\,
            sr => \N__49519\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__40341\,
            in1 => \N__40464\,
            in2 => \_gnd_net_\,
            in3 => \N__40345\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => \N__40327\,
            sr => \N__49519\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__40264\,
            in1 => \N__44785\,
            in2 => \N__41031\,
            in3 => \N__40778\,
            lcout => \elapsed_time_ns_1_RNI3JIF91_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__44416\,
            in1 => \N__40285\,
            in2 => \N__41029\,
            in3 => \N__40776\,
            lcout => \elapsed_time_ns_1_RNIQ9IF91_0_20\,
            ltout => \elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40278\,
            in1 => \N__40563\,
            in2 => \N__40267\,
            in3 => \N__40263\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__44293\,
            in1 => \N__40249\,
            in2 => \N__41030\,
            in3 => \N__40777\,
            lcout => \elapsed_time_ns_1_RNITCIF91_0_23\,
            ltout => \elapsed_time_ns_1_RNITCIF91_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40584\,
            in2 => \N__40600\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__41033\,
            in1 => \N__44248\,
            in2 => \N__40588\,
            in3 => \N__40783\,
            lcout => \elapsed_time_ns_1_RNIUDIF91_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__43929\,
            in1 => \N__47152\,
            in2 => \N__47776\,
            in3 => \N__40705\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010001"
        )
    port map (
            in0 => \N__44680\,
            in1 => \N__40861\,
            in2 => \N__40573\,
            in3 => \N__40839\,
            lcout => \delay_measurement_inst.delay_tr9\,
            ltout => \delay_measurement_inst.delay_tr9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__47743\,
            in1 => \N__40638\,
            in2 => \N__40570\,
            in3 => \N__41034\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__41035\,
            in1 => \N__41443\,
            in2 => \N__45334\,
            in3 => \N__47775\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__40782\,
            in1 => \N__41032\,
            in2 => \N__40567\,
            in3 => \N__44722\,
            lcout => \elapsed_time_ns_1_RNIRBJF91_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__41039\,
            in1 => \N__41488\,
            in2 => \N__45332\,
            in3 => \N__47233\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__41318\,
            in1 => \N__47794\,
            in2 => \N__45335\,
            in3 => \N__41042\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__41040\,
            in1 => \N__41096\,
            in2 => \N__47410\,
            in3 => \N__40787\,
            lcout => \elapsed_time_ns_1_RNICG2591_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJL0B1_24_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__44721\,
            in1 => \N__44784\,
            in2 => \_gnd_net_\,
            in3 => \N__44244\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_23_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44289\,
            in1 => \N__44157\,
            in2 => \N__40843\,
            in3 => \N__40870\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__40786\,
            in1 => \N__47422\,
            in2 => \N__41139\,
            in3 => \N__41041\,
            lcout => \elapsed_time_ns_1_RNIDH2591_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__47793\,
            in1 => \N__40606\,
            in2 => \_gnd_net_\,
            in3 => \N__47245\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__47212\,
            in1 => \N__41963\,
            in2 => \N__45336\,
            in3 => \N__41043\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101110"
        )
    port map (
            in0 => \N__40684\,
            in1 => \N__41361\,
            in2 => \N__47386\,
            in3 => \N__41045\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40699\,
            in3 => \N__45333\,
            lcout => \elapsed_time_ns_1_RNIK8NQL1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__40651\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41359\,
            lcout => \elapsed_time_ns_1_RNINBNQL1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44094\,
            in1 => \N__44046\,
            in2 => \N__44007\,
            in3 => \N__43476\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_353\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_353_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43916\,
            in1 => \N__47292\,
            in2 => \N__41176\,
            in3 => \N__47265\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__41360\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41155\,
            lcout => \elapsed_time_ns_1_RNI8765M1_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41358\,
            in2 => \_gnd_net_\,
            in3 => \N__41149\,
            lcout => \elapsed_time_ns_1_RNIA965M1_0_18\,
            ltout => \elapsed_time_ns_1_RNIA965M1_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41860\,
            in1 => \N__41125\,
            in2 => \N__41107\,
            in3 => \N__41089\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40888\,
            in2 => \_gnd_net_\,
            in3 => \N__41362\,
            lcout => \elapsed_time_ns_1_RNI9865M1_0_17\,
            ltout => \elapsed_time_ns_1_RNI9865M1_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__47193\,
            in1 => \N__41044\,
            in2 => \N__40891\,
            in3 => \N__45314\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40882\,
            in2 => \_gnd_net_\,
            in3 => \N__41364\,
            lcout => \elapsed_time_ns_1_RNIBA65M1_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG7AP1_20_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44907\,
            in1 => \N__44196\,
            in2 => \N__44853\,
            in3 => \N__44409\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__44331\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44370\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lt31_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__41363\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41458\,
            lcout => \elapsed_time_ns_1_RNI6565M1_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__49582\,
            in1 => \N__41391\,
            in2 => \N__44692\,
            in3 => \N__41376\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__41332\,
            in1 => \_gnd_net_\,
            in2 => \N__41323\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIQENQL1_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__50292\,
            in1 => \N__45184\,
            in2 => \N__50038\,
            in3 => \N__47679\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41262\,
            in2 => \_gnd_net_\,
            in3 => \N__41222\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_hc_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__44552\,
            in1 => \N__41274\,
            in2 => \N__41281\,
            in3 => \N__46152\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46135\,
            in2 => \_gnd_net_\,
            in3 => \N__46151\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_RNIG7JF_2_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41189\,
            in2 => \_gnd_net_\,
            in3 => \N__46190\,
            lcout => \phase_controller_inst2.state_RNIG7JFZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_2_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__41190\,
            in1 => \N__41263\,
            in2 => \N__46197\,
            in3 => \N__41223\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49434\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__47814\,
            in1 => \N__48093\,
            in2 => \N__41887\,
            in3 => \N__41932\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__41931\,
            in1 => \N__47815\,
            in2 => \N__48097\,
            in3 => \N__41883\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001000110010"
        )
    port map (
            in0 => \N__41967\,
            in1 => \N__41798\,
            in2 => \N__41655\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49922\,
            ce => \N__50320\,
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__41799\,
            in1 => \N__41922\,
            in2 => \_gnd_net_\,
            in3 => \N__41647\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49922\,
            ce => \N__50320\,
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001000110010"
        )
    port map (
            in0 => \N__41868\,
            in1 => \N__41801\,
            in2 => \N__41656\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49922\,
            ce => \N__50320\,
            sr => \N__49440\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100001101"
        )
    port map (
            in0 => \N__48069\,
            in1 => \N__41467\,
            in2 => \N__48046\,
            in3 => \N__41823\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__41466\,
            in1 => \N__48042\,
            in2 => \N__41827\,
            in3 => \N__48070\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__41800\,
            in1 => \N__41648\,
            in2 => \_gnd_net_\,
            in3 => \N__41502\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49922\,
            ce => \N__50320\,
            sr => \N__49440\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__42382\,
            in1 => \N__45903\,
            in2 => \N__43259\,
            in3 => \N__45466\,
            lcout => \elapsed_time_ns_1_RNI3ET8E1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__45311\,
            in1 => \N__49584\,
            in2 => \_gnd_net_\,
            in3 => \N__42363\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__42400\,
            in1 => \N__43208\,
            in2 => \N__42100\,
            in3 => \N__45465\,
            lcout => \elapsed_time_ns_1_RNI4FT8E1_0_12\,
            ltout => \elapsed_time_ns_1_RNI4FT8E1_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44971\,
            in1 => \N__43249\,
            in2 => \N__42097\,
            in3 => \N__43298\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42094\,
            in1 => \N__42082\,
            in2 => \N__42070\,
            in3 => \N__45043\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__44664\,
            in1 => \N__42135\,
            in2 => \N__42055\,
            in3 => \N__47718\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_369\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42052\,
            in3 => \N__45312\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_367_clk\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_367_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__45902\,
            in1 => \N__42015\,
            in2 => \N__42049\,
            in3 => \N__42046\,
            lcout => \elapsed_time_ns_1_RNI3FU8E1_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42345\,
            in1 => \N__42033\,
            in2 => \N__42016\,
            in3 => \N__42117\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__45463\,
            in1 => \N__42346\,
            in2 => \N__42454\,
            in3 => \N__45874\,
            lcout => \elapsed_time_ns_1_RNI5HU8E1_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__45872\,
            in1 => \N__45462\,
            in2 => \N__42421\,
            in3 => \N__45123\,
            lcout => \elapsed_time_ns_1_RNI6IU8E1_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__45461\,
            in1 => \N__45148\,
            in2 => \N__42436\,
            in3 => \N__45873\,
            lcout => \elapsed_time_ns_1_RNI7JU8E1_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__42306\,
            in1 => \N__45460\,
            in2 => \N__45906\,
            in3 => \N__42327\,
            lcout => \elapsed_time_ns_1_RNIMHKEE1_0_5\,
            ltout => \elapsed_time_ns_1_RNIMHKEE1_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__47076\,
            in1 => \N__42286\,
            in2 => \N__42223\,
            in3 => \N__42216\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49911\,
            ce => \N__48951\,
            sr => \N__49458\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__42136\,
            in1 => \N__47077\,
            in2 => \N__45907\,
            in3 => \N__45464\,
            lcout => \elapsed_time_ns_1_RNI5IV8E1_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__42962\,
            in1 => \N__42118\,
            in2 => \N__45353\,
            in3 => \N__45514\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42103\,
            in3 => \N__46000\,
            lcout => \elapsed_time_ns_1_RNIIIC6P1_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__45096\,
            in1 => \N__42496\,
            in2 => \N__45549\,
            in3 => \N__45915\,
            lcout => \elapsed_time_ns_1_RNI9LU8E1_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__45513\,
            in1 => \N__42546\,
            in2 => \N__45928\,
            in3 => \N__42487\,
            lcout => \elapsed_time_ns_1_RNIBNU8E1_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__42526\,
            in1 => \N__45911\,
            in2 => \N__42505\,
            in3 => \N__45512\,
            lcout => \elapsed_time_ns_1_RNIAMU8E1_0_27\,
            ltout => \elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42495\,
            in1 => \N__42486\,
            in2 => \N__42478\,
            in3 => \N__42471\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42460\,
            in1 => \N__42450\,
            in2 => \N__42439\,
            in3 => \N__42406\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42432\,
            in2 => \_gnd_net_\,
            in3 => \N__42417\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45006\,
            in1 => \N__42399\,
            in2 => \N__42592\,
            in3 => \N__42378\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__42367\,
            in1 => \N__49585\,
            in2 => \_gnd_net_\,
            in3 => \N__45313\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_344_i\,
            ltout => \delay_measurement_inst.delay_hc_timer.N_344_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42352\,
            in3 => \N__42598\,
            lcout => \elapsed_time_ns_1_RNIHHC6P1_0_18\,
            ltout => \elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__42955\,
            in1 => \N__42773\,
            in2 => \N__42349\,
            in3 => \N__42643\,
            lcout => \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42789\,
            in1 => \N__45801\,
            in2 => \N__42610\,
            in3 => \N__42573\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010111010"
        )
    port map (
            in0 => \N__45315\,
            in1 => \N__45524\,
            in2 => \N__43376\,
            in3 => \N__42609\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101100"
        )
    port map (
            in0 => \N__42591\,
            in1 => \N__45316\,
            in2 => \N__45550\,
            in3 => \N__46884\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42580\,
            in3 => \N__46013\,
            lcout => \elapsed_time_ns_1_RNIDDC6P1_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__42644\,
            in1 => \N__45545\,
            in2 => \N__45352\,
            in3 => \N__42577\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42562\,
            in3 => \N__46004\,
            lcout => \elapsed_time_ns_1_RNIFFC6P1_0_16\,
            ltout => \elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46794\,
            in2 => \N__42559\,
            in3 => \N__47055\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49897\,
            ce => \N__49108\,
            sr => \N__49482\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__42555\,
            in1 => \N__48495\,
            in2 => \N__48523\,
            in3 => \N__42801\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__48496\,
            in1 => \N__48519\,
            in2 => \N__42805\,
            in3 => \N__42556\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__47056\,
            in1 => \_gnd_net_\,
            in2 => \N__46827\,
            in3 => \N__42774\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49897\,
            ce => \N__49108\,
            sr => \N__49482\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__42964\,
            in1 => \N__47057\,
            in2 => \_gnd_net_\,
            in3 => \N__46795\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49897\,
            ce => \N__49108\,
            sr => \N__49482\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__42928\,
            in1 => \N__48665\,
            in2 => \N__48475\,
            in3 => \N__42909\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__42769\,
            in1 => \N__45546\,
            in2 => \N__45364\,
            in3 => \N__42793\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42778\,
            in3 => \N__46016\,
            lcout => \elapsed_time_ns_1_RNIGGC6P1_0_17\,
            ltout => \elapsed_time_ns_1_RNIGGC6P1_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__47059\,
            in1 => \_gnd_net_\,
            in2 => \N__42742\,
            in3 => \N__46810\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49891\,
            ce => \N__43148\,
            sr => \N__49489\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__42681\,
            in1 => \N__42618\,
            in2 => \N__42721\,
            in3 => \N__42690\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__42619\,
            in1 => \N__42717\,
            in2 => \N__42694\,
            in3 => \N__42682\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__42645\,
            in1 => \N__47058\,
            in2 => \_gnd_net_\,
            in3 => \N__46799\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49891\,
            ce => \N__43148\,
            sr => \N__49489\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__47060\,
            in1 => \N__46811\,
            in2 => \_gnd_net_\,
            in3 => \N__42963\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49891\,
            ce => \N__43148\,
            sr => \N__49489\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__45735\,
            in1 => \N__46885\,
            in2 => \_gnd_net_\,
            in3 => \N__45673\,
            lcout => \phase_controller_inst1.stoper_hc.N_318\,
            ltout => \phase_controller_inst1.stoper_hc.N_318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__47062\,
            in1 => \N__43308\,
            in2 => \N__42931\,
            in3 => \N__46806\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49883\,
            ce => \N__49123\,
            sr => \N__49494\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__46802\,
            in1 => \N__47063\,
            in2 => \N__43264\,
            in3 => \N__46922\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49883\,
            ce => \N__49123\,
            sr => \N__49494\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__47064\,
            in1 => \N__46805\,
            in2 => \N__46930\,
            in3 => \N__43215\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49883\,
            ce => \N__49123\,
            sr => \N__49494\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__46803\,
            in1 => \N__47065\,
            in2 => \N__44995\,
            in3 => \N__46923\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49883\,
            ce => \N__49123\,
            sr => \N__49494\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010001010100"
        )
    port map (
            in0 => \N__47061\,
            in1 => \N__46804\,
            in2 => \N__43381\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49883\,
            ce => \N__49123\,
            sr => \N__49494\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000100"
        )
    port map (
            in0 => \N__48474\,
            in1 => \N__42927\,
            in2 => \N__48673\,
            in3 => \N__42913\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010110010"
        )
    port map (
            in0 => \N__42894\,
            in1 => \N__42874\,
            in2 => \N__43344\,
            in3 => \N__42850\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__47066\,
            in1 => \N__46822\,
            in2 => \_gnd_net_\,
            in3 => \N__43377\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => \N__43149\,
            sr => \N__49504\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__46926\,
            in1 => \N__47072\,
            in2 => \N__46831\,
            in3 => \N__46890\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => \N__43149\,
            sr => \N__49504\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__47068\,
            in1 => \N__46927\,
            in2 => \N__43309\,
            in3 => \N__46825\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => \N__43149\,
            sr => \N__49504\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__46924\,
            in1 => \N__47069\,
            in2 => \N__46829\,
            in3 => \N__43263\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => \N__43149\,
            sr => \N__49504\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__47070\,
            in1 => \N__46823\,
            in2 => \N__43219\,
            in3 => \N__46928\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => \N__43149\,
            sr => \N__49504\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__46925\,
            in1 => \N__47071\,
            in2 => \N__46830\,
            in3 => \N__44994\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => \N__43149\,
            sr => \N__49504\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__47067\,
            in1 => \N__45756\,
            in2 => \N__45610\,
            in3 => \N__46824\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49877\,
            ce => \N__43149\,
            sr => \N__49504\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43822\,
            in1 => \N__46520\,
            in2 => \_gnd_net_\,
            in3 => \N__42970\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__49966\,
            ce => \N__43687\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43818\,
            in1 => \N__47498\,
            in2 => \_gnd_net_\,
            in3 => \N__42967\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__49966\,
            ce => \N__43687\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43823\,
            in1 => \N__43620\,
            in2 => \_gnd_net_\,
            in3 => \N__43408\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__49966\,
            ce => \N__43687\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43819\,
            in1 => \N__43596\,
            in2 => \_gnd_net_\,
            in3 => \N__43405\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__49966\,
            ce => \N__43687\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43824\,
            in1 => \N__43571\,
            in2 => \_gnd_net_\,
            in3 => \N__43402\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__49966\,
            ce => \N__43687\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43820\,
            in1 => \N__43544\,
            in2 => \_gnd_net_\,
            in3 => \N__43399\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__49966\,
            ce => \N__43687\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43825\,
            in1 => \N__43518\,
            in2 => \_gnd_net_\,
            in3 => \N__43396\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__49966\,
            ce => \N__43687\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43821\,
            in1 => \N__43494\,
            in2 => \_gnd_net_\,
            in3 => \N__43393\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__49966\,
            ce => \N__43687\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43772\,
            in1 => \N__44120\,
            in2 => \_gnd_net_\,
            in3 => \N__43390\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__49961\,
            ce => \N__43683\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43776\,
            in1 => \N__44072\,
            in2 => \_gnd_net_\,
            in3 => \N__43387\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__49961\,
            ce => \N__43683\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43769\,
            in1 => \N__44025\,
            in2 => \_gnd_net_\,
            in3 => \N__43384\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__49961\,
            ce => \N__43683\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43773\,
            in1 => \N__43973\,
            in2 => \_gnd_net_\,
            in3 => \N__43435\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__49961\,
            ce => \N__43683\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43770\,
            in1 => \N__43946\,
            in2 => \_gnd_net_\,
            in3 => \N__43432\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__49961\,
            ce => \N__43683\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43774\,
            in1 => \N__43898\,
            in2 => \_gnd_net_\,
            in3 => \N__43429\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__49961\,
            ce => \N__43683\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43771\,
            in1 => \N__43872\,
            in2 => \_gnd_net_\,
            in3 => \N__43426\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__49961\,
            ce => \N__43683\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43775\,
            in1 => \N__43842\,
            in2 => \_gnd_net_\,
            in3 => \N__43423\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__49961\,
            ce => \N__43683\,
            sr => \N__49409\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43777\,
            in1 => \N__44462\,
            in2 => \_gnd_net_\,
            in3 => \N__43420\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__49955\,
            ce => \N__43676\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43814\,
            in1 => \N__44435\,
            in2 => \_gnd_net_\,
            in3 => \N__43417\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__49955\,
            ce => \N__43676\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43778\,
            in1 => \N__44393\,
            in2 => \_gnd_net_\,
            in3 => \N__43414\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__49955\,
            ce => \N__43676\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43815\,
            in1 => \N__44354\,
            in2 => \_gnd_net_\,
            in3 => \N__43411\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__49955\,
            ce => \N__43676\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43779\,
            in1 => \N__44309\,
            in2 => \_gnd_net_\,
            in3 => \N__43462\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__49955\,
            ce => \N__43676\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43816\,
            in1 => \N__44264\,
            in2 => \_gnd_net_\,
            in3 => \N__43459\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__49955\,
            ce => \N__43676\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43780\,
            in1 => \N__44220\,
            in2 => \_gnd_net_\,
            in3 => \N__43456\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__49955\,
            ce => \N__43676\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43817\,
            in1 => \N__44175\,
            in2 => \_gnd_net_\,
            in3 => \N__43453\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__49955\,
            ce => \N__43676\,
            sr => \N__49411\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43808\,
            in1 => \N__44933\,
            in2 => \_gnd_net_\,
            in3 => \N__43450\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__49950\,
            ce => \N__43675\,
            sr => \N__49413\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43812\,
            in1 => \N__44876\,
            in2 => \_gnd_net_\,
            in3 => \N__43447\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__49950\,
            ce => \N__43675\,
            sr => \N__49413\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43809\,
            in1 => \N__44804\,
            in2 => \_gnd_net_\,
            in3 => \N__43444\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__49950\,
            ce => \N__43675\,
            sr => \N__49413\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43813\,
            in1 => \N__44758\,
            in2 => \_gnd_net_\,
            in3 => \N__43441\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__49950\,
            ce => \N__43675\,
            sr => \N__49413\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43810\,
            in1 => \N__44823\,
            in2 => \_gnd_net_\,
            in3 => \N__43438\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__49950\,
            ce => \N__43675\,
            sr => \N__49413\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__44736\,
            in1 => \N__43811\,
            in2 => \_gnd_net_\,
            in3 => \N__43690\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49950\,
            ce => \N__43675\,
            sr => \N__49413\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43626\,
            in2 => \N__46534\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49946\,
            ce => \N__47475\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43602\,
            in2 => \N__47512\,
            in3 => \N__43630\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49946\,
            ce => \N__47475\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43627\,
            in2 => \N__43578\,
            in3 => \N__43606\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49946\,
            ce => \N__47475\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43603\,
            in2 => \N__43551\,
            in3 => \N__43582\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49946\,
            ce => \N__47475\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43524\,
            in2 => \N__43579\,
            in3 => \N__43555\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49946\,
            ce => \N__47475\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43500\,
            in2 => \N__43552\,
            in3 => \N__43528\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49946\,
            ce => \N__47475\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43525\,
            in2 => \N__44127\,
            in3 => \N__43504\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49946\,
            ce => \N__47475\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43501\,
            in2 => \N__44079\,
            in3 => \N__43465\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49946\,
            ce => \N__47475\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44031\,
            in2 => \N__44131\,
            in3 => \N__44083\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49941\,
            ce => \N__47477\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43980\,
            in2 => \N__44080\,
            in3 => \N__44035\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49941\,
            ce => \N__47477\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44032\,
            in2 => \N__43953\,
            in3 => \N__43990\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49941\,
            ce => \N__47477\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43899\,
            in2 => \N__43987\,
            in3 => \N__43957\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49941\,
            ce => \N__47477\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43878\,
            in2 => \N__43954\,
            in3 => \N__43903\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr9lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49941\,
            ce => \N__47477\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43900\,
            in2 => \N__43854\,
            in3 => \N__43882\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49941\,
            ce => \N__47477\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43879\,
            in2 => \N__44475\,
            in3 => \N__43858\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49941\,
            ce => \N__47477\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44436\,
            in2 => \N__43855\,
            in3 => \N__43828\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49941\,
            ce => \N__47477\,
            sr => \N__49423\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44394\,
            in2 => \N__44476\,
            in3 => \N__44446\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49934\,
            ce => \N__47478\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44355\,
            in2 => \N__44443\,
            in3 => \N__44398\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49934\,
            ce => \N__47478\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44395\,
            in2 => \N__44316\,
            in3 => \N__44359\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49934\,
            ce => \N__47478\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44356\,
            in2 => \N__44271\,
            in3 => \N__44320\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49934\,
            ce => \N__47478\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44226\,
            in2 => \N__44317\,
            in3 => \N__44275\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49934\,
            ce => \N__47478\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44181\,
            in2 => \N__44272\,
            in3 => \N__44230\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49934\,
            ce => \N__47478\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44227\,
            in2 => \N__44940\,
            in3 => \N__44185\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49934\,
            ce => \N__47478\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44182\,
            in2 => \N__44883\,
            in3 => \N__44134\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49934\,
            ce => \N__47478\,
            sr => \N__49425\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44805\,
            in2 => \N__44941\,
            in3 => \N__44890\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49929\,
            ce => \N__47479\,
            sr => \N__49435\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44756\,
            in2 => \N__44887\,
            in3 => \N__44827\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49929\,
            ce => \N__47479\,
            sr => \N__49435\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44824\,
            in2 => \N__44809\,
            in3 => \N__44761\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49929\,
            ce => \N__47479\,
            sr => \N__49435\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44757\,
            in2 => \N__44740\,
            in3 => \N__44701\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49929\,
            ce => \N__47479\,
            sr => \N__49435\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44698\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49929\,
            ce => \N__47479\,
            sr => \N__49435\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__44641\,
            in1 => \N__46665\,
            in2 => \N__46606\,
            in3 => \N__44597\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__44557\,
            in1 => \N__44503\,
            in2 => \N__44479\,
            in3 => \N__50131\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49923\,
            ce => 'H',
            sr => \N__49441\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110101"
        )
    port map (
            in0 => \N__50106\,
            in1 => \N__48200\,
            in2 => \N__48171\,
            in3 => \N__45196\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45187\,
            in3 => \N__50017\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50018\,
            in2 => \_gnd_net_\,
            in3 => \N__45180\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45168\,
            in1 => \N__45147\,
            in2 => \N__45127\,
            in3 => \N__45097\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__45076\,
            in1 => \N__45070\,
            in2 => \N__45058\,
            in3 => \N__45055\,
            lcout => \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__48231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48216\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__48261\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48246\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__45013\,
            in1 => \N__45922\,
            in2 => \N__44987\,
            in3 => \N__45470\,
            lcout => \elapsed_time_ns_1_RNI5GT8E1_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48166\,
            in2 => \_gnd_net_\,
            in3 => \N__48201\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__45374\,
            in1 => \N__45958\,
            in2 => \N__45552\,
            in3 => \N__46047\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46027\,
            in3 => \N__46014\,
            lcout => \elapsed_time_ns_1_RNIUE3CP1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__45701\,
            in1 => \N__45926\,
            in2 => \N__45551\,
            in3 => \N__45808\,
            lcout => \elapsed_time_ns_1_RNI7IT8E1_0_15\,
            ltout => \elapsed_time_ns_1_RNI7IT8E1_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.N_269_i_1_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010100"
        )
    port map (
            in0 => \N__45654\,
            in1 => \N__46870\,
            in2 => \N__45790\,
            in3 => \N__45779\,
            lcout => \phase_controller_inst1.stoper_hc.N_269_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__47020\,
            in1 => \N__46745\,
            in2 => \N__45717\,
            in3 => \N__45655\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => \N__48993\,
            sr => \N__49459\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__45630\,
            in1 => \N__45609\,
            in2 => \N__45556\,
            in3 => \N__45375\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46218\,
            in2 => \_gnd_net_\,
            in3 => \N__46245\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110101"
        )
    port map (
            in0 => \N__46126\,
            in1 => \N__48736\,
            in2 => \N__48715\,
            in3 => \N__47140\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46252\,
            in3 => \N__46219\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__46220\,
            in1 => \N__48994\,
            in2 => \N__46249\,
            in3 => \N__48142\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49465\
        );

    \phase_controller_inst2.stoper_hc.running_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001111110000"
        )
    port map (
            in0 => \N__47124\,
            in1 => \N__46127\,
            in2 => \N__46237\,
            in3 => \N__46221\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49465\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__46125\,
            in1 => \N__46233\,
            in2 => \_gnd_net_\,
            in3 => \N__46158\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110000001100"
        )
    port map (
            in0 => \N__47125\,
            in1 => \N__46181\,
            in2 => \N__46225\,
            in3 => \N__46128\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49465\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46159\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49465\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46108\,
            in2 => \N__46099\,
            in3 => \N__48140\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46090\,
            in2 => \N__46078\,
            in3 => \N__48115\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48435\,
            in1 => \N__46069\,
            in2 => \N__46057\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46411\,
            in2 => \N__46402\,
            in3 => \N__48415\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46393\,
            in2 => \N__46381\,
            in3 => \N__48397\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48379\,
            in1 => \N__46369\,
            in2 => \N__46354\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46345\,
            in2 => \N__46330\,
            in3 => \N__48361\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48343\,
            in1 => \N__46318\,
            in2 => \N__46309\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48325\,
            in1 => \N__46300\,
            in2 => \N__46291\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46282\,
            in2 => \N__46276\,
            in3 => \N__48307\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48616\,
            in1 => \N__46267\,
            in2 => \N__46261\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46492\,
            in2 => \N__46501\,
            in3 => \N__48595\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46486\,
            in2 => \N__46480\,
            in3 => \N__48577\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48559\,
            in1 => \N__46471\,
            in2 => \N__46678\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46465\,
            in2 => \N__46456\,
            in3 => \N__48541\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46447\,
            in2 => \N__46441\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46429\,
            in2 => \N__46420\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50329\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48772\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50365\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48808\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48742\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48679\,
            in2 => \N__48711\,
            in3 => \N__47131\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47128\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__47113\,
            in1 => \N__46929\,
            in2 => \N__46891\,
            in3 => \N__46828\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49884\,
            ce => \N__49069\,
            sr => \N__49495\
        );

    \phase_controller_inst1.T12_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__46545\,
            in1 => \N__46666\,
            in2 => \_gnd_net_\,
            in3 => \N__46599\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49878\,
            ce => 'H',
            sr => \N__49505\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46533\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => \N__47476\,
            sr => \N__49412\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47511\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => \N__47476\,
            sr => \N__49412\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__47382\,
            in1 => \N__47762\,
            in2 => \N__47364\,
            in3 => \N__47791\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_19_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__47172\,
            in1 => \N__47428\,
            in2 => \N__47458\,
            in3 => \N__47395\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2BNE1_16_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47226\,
            in1 => \N__47189\,
            in2 => \N__47742\,
            in3 => \N__47207\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47421\,
            in2 => \_gnd_net_\,
            in3 => \N__47406\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_346\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47381\,
            in1 => \N__47351\,
            in2 => \N__47335\,
            in3 => \N__47322\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_349\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_349_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__47291\,
            in1 => \N__47264\,
            in2 => \N__47248\,
            in3 => \N__47734\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__47225\,
            in1 => \N__47208\,
            in2 => \N__47194\,
            in3 => \N__47171\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_362\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__47792\,
            in1 => \N__47763\,
            in2 => \N__47746\,
            in3 => \N__47738\,
            lcout => \delay_measurement_inst.N_365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47689\,
            in2 => \N__47680\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50288\,
            in1 => \N__47655\,
            in2 => \_gnd_net_\,
            in3 => \N__47641\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__50293\,
            in1 => \N__47622\,
            in2 => \N__47638\,
            in3 => \N__47608\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50289\,
            in1 => \N__47601\,
            in2 => \_gnd_net_\,
            in3 => \N__47587\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50294\,
            in1 => \N__47583\,
            in2 => \_gnd_net_\,
            in3 => \N__47569\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50290\,
            in1 => \N__47565\,
            in2 => \_gnd_net_\,
            in3 => \N__47551\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50295\,
            in1 => \N__47544\,
            in2 => \_gnd_net_\,
            in3 => \N__47530\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50291\,
            in1 => \N__47526\,
            in2 => \_gnd_net_\,
            in3 => \N__47944\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49424\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50276\,
            in1 => \N__47940\,
            in2 => \_gnd_net_\,
            in3 => \N__47926\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50269\,
            in1 => \N__47922\,
            in2 => \_gnd_net_\,
            in3 => \N__47908\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50273\,
            in1 => \N__47904\,
            in2 => \_gnd_net_\,
            in3 => \N__47890\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50270\,
            in1 => \N__47886\,
            in2 => \_gnd_net_\,
            in3 => \N__47872\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50274\,
            in1 => \N__47868\,
            in2 => \_gnd_net_\,
            in3 => \N__47854\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50271\,
            in1 => \N__47850\,
            in2 => \_gnd_net_\,
            in3 => \N__47836\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50275\,
            in1 => \N__47832\,
            in2 => \_gnd_net_\,
            in3 => \N__47818\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50272\,
            in1 => \N__47813\,
            in2 => \_gnd_net_\,
            in3 => \N__47797\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49426\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50277\,
            in1 => \N__48087\,
            in2 => \_gnd_net_\,
            in3 => \N__48073\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50281\,
            in1 => \N__48063\,
            in2 => \_gnd_net_\,
            in3 => \N__48049\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50278\,
            in1 => \N__48036\,
            in2 => \_gnd_net_\,
            in3 => \N__48022\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50282\,
            in1 => \N__48861\,
            in2 => \_gnd_net_\,
            in3 => \N__48019\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50279\,
            in1 => \N__48876\,
            in2 => \_gnd_net_\,
            in3 => \N__48016\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50283\,
            in1 => \N__48009\,
            in2 => \_gnd_net_\,
            in3 => \N__47995\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50280\,
            in1 => \N__47985\,
            in2 => \_gnd_net_\,
            in3 => \N__47971\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50284\,
            in1 => \N__47961\,
            in2 => \_gnd_net_\,
            in3 => \N__47947\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49436\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50301\,
            in1 => \N__48279\,
            in2 => \_gnd_net_\,
            in3 => \N__48265\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49442\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50305\,
            in1 => \N__48262\,
            in2 => \_gnd_net_\,
            in3 => \N__48250\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49442\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50302\,
            in1 => \N__48247\,
            in2 => \_gnd_net_\,
            in3 => \N__48235\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49442\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50306\,
            in1 => \N__48232\,
            in2 => \_gnd_net_\,
            in3 => \N__48220\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49442\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50303\,
            in1 => \N__48217\,
            in2 => \_gnd_net_\,
            in3 => \N__48205\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49442\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50307\,
            in1 => \N__48202\,
            in2 => \_gnd_net_\,
            in3 => \N__48184\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49442\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50304\,
            in1 => \N__48170\,
            in2 => \_gnd_net_\,
            in3 => \N__48181\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49442\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48141\,
            in2 => \N__48124\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48983\,
            in1 => \N__48114\,
            in2 => \_gnd_net_\,
            in3 => \N__48100\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__48961\,
            in1 => \N__48442\,
            in2 => \N__48436\,
            in3 => \N__48418\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48984\,
            in1 => \N__48414\,
            in2 => \_gnd_net_\,
            in3 => \N__48400\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48962\,
            in1 => \N__48396\,
            in2 => \_gnd_net_\,
            in3 => \N__48382\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48985\,
            in1 => \N__48378\,
            in2 => \_gnd_net_\,
            in3 => \N__48364\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48963\,
            in1 => \N__48360\,
            in2 => \_gnd_net_\,
            in3 => \N__48346\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48986\,
            in1 => \N__48342\,
            in2 => \_gnd_net_\,
            in3 => \N__48328\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49451\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49104\,
            in1 => \N__48324\,
            in2 => \_gnd_net_\,
            in3 => \N__48310\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49079\,
            in1 => \N__48303\,
            in2 => \_gnd_net_\,
            in3 => \N__48289\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49101\,
            in1 => \N__48615\,
            in2 => \_gnd_net_\,
            in3 => \N__48598\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49080\,
            in1 => \N__48594\,
            in2 => \_gnd_net_\,
            in3 => \N__48580\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49102\,
            in1 => \N__48576\,
            in2 => \_gnd_net_\,
            in3 => \N__48562\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49081\,
            in1 => \N__48558\,
            in2 => \_gnd_net_\,
            in3 => \N__48544\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49103\,
            in1 => \N__48540\,
            in2 => \_gnd_net_\,
            in3 => \N__48526\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49082\,
            in1 => \N__48513\,
            in2 => \_gnd_net_\,
            in3 => \N__48499\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49460\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49083\,
            in1 => \N__48494\,
            in2 => \_gnd_net_\,
            in3 => \N__48478\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49087\,
            in1 => \N__48467\,
            in2 => \_gnd_net_\,
            in3 => \N__48445\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49084\,
            in1 => \N__48669\,
            in2 => \_gnd_net_\,
            in3 => \N__48643\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49088\,
            in1 => \N__50343\,
            in2 => \_gnd_net_\,
            in3 => \N__48640\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49085\,
            in1 => \N__50358\,
            in2 => \_gnd_net_\,
            in3 => \N__48637\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49089\,
            in1 => \N__48786\,
            in2 => \_gnd_net_\,
            in3 => \N__48634\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49086\,
            in1 => \N__48801\,
            in2 => \_gnd_net_\,
            in3 => \N__48631\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49090\,
            in1 => \N__50379\,
            in2 => \_gnd_net_\,
            in3 => \N__48628\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49908\,
            ce => 'H',
            sr => \N__49466\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49098\,
            in1 => \N__50392\,
            in2 => \_gnd_net_\,
            in3 => \N__48625\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49091\,
            in1 => \N__48820\,
            in2 => \_gnd_net_\,
            in3 => \N__48622\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49099\,
            in1 => \N__48832\,
            in2 => \_gnd_net_\,
            in3 => \N__48619\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49092\,
            in1 => \N__48754\,
            in2 => \_gnd_net_\,
            in3 => \N__49132\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49100\,
            in1 => \N__48766\,
            in2 => \_gnd_net_\,
            in3 => \N__49129\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__49093\,
            in1 => \N__48735\,
            in2 => \_gnd_net_\,
            in3 => \N__49126\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49473\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__48706\,
            in1 => \N__49094\,
            in2 => \_gnd_net_\,
            in3 => \N__48883\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49473\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48880\,
            in2 => \_gnd_net_\,
            in3 => \N__48862\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48831\,
            in2 => \_gnd_net_\,
            in3 => \N__48819\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48802\,
            in2 => \_gnd_net_\,
            in3 => \N__48787\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48765\,
            in2 => \_gnd_net_\,
            in3 => \N__48753\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__48734\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48710\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50391\,
            in2 => \_gnd_net_\,
            in3 => \N__50380\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50359\,
            in2 => \_gnd_net_\,
            in3 => \N__50344\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_df20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50102\,
            in2 => \_gnd_net_\,
            in3 => \N__50139\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__50088\,
            in1 => \N__49989\,
            in2 => \_gnd_net_\,
            in3 => \N__50132\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50140\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49936\,
            ce => 'H',
            sr => \N__49443\
        );

    \phase_controller_inst1.stoper_tr.running_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__50098\,
            in1 => \N__50062\,
            in2 => \N__49993\,
            in3 => \N__50016\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49936\,
            ce => 'H',
            sr => \N__49443\
        );
end \INTERFACE\;
